/* rom.v : rom */

module rom
#(parameter BITS = 16, ADDRESS_BITS = 8)
(
	input CLK,
	input [ADDRESS_BITS - 1 : 0]  ADDRESS,
	output [BITS - 1 : 0] DATA_OUT,
);

localparam ROM_ADDRESS_BITS = 8;

reg [BITS - 1:0] mem [(1 << ROM_ADDRESS_BITS) - 1:0];
reg [BITS - 1:0] dout;
assign DATA_OUT = dout;
initial mem[0] = 16'h1002;
initial mem[1] = 16'h4600;
initial mem[2] = 16'h1007;
initial mem[3] = 16'h4608;
initial mem[4] = 16'h1007;
initial mem[5] = 16'h4608;
initial mem[6] = 16'h1007;
initial mem[7] = 16'h4608;
initial mem[8] = 16'h1007;
initial mem[9] = 16'h4608;
initial mem[10] = 16'h0000;
initial mem[11] = 16'h0000;
initial mem[12] = 16'h0000;
initial mem[13] = 16'h0000;
initial mem[14] = 16'h0000;
initial mem[15] = 16'h0000;
initial mem[16] = 16'h0000;
initial mem[17] = 16'h0000;
initial mem[18] = 16'h0000;
initial mem[19] = 16'h0000;
initial mem[20] = 16'h0000;
initial mem[21] = 16'h0000;
initial mem[22] = 16'h0000;
initial mem[23] = 16'h0000;
initial mem[24] = 16'h0000;
initial mem[25] = 16'h0000;
initial mem[26] = 16'h0000;
initial mem[27] = 16'h0000;
initial mem[28] = 16'h0000;
initial mem[29] = 16'h0000;
initial mem[30] = 16'h0000;
initial mem[31] = 16'h0000;
initial mem[32] = 16'h1003;
initial mem[33] = 16'h301b;
initial mem[34] = 16'h1000;
initial mem[35] = 16'h3028;
initial mem[36] = 16'h2060;
initial mem[37] = 16'hc230;
initial mem[38] = 16'h3111;
initial mem[39] = 16'h1540;
initial mem[40] = 16'hed30;
initial mem[41] = 16'h3161;
initial mem[42] = 16'h3321;
initial mem[43] = 16'h1002;
initial mem[44] = 16'h4105;
initial mem[45] = 16'h3041;
initial mem[46] = 16'h15d2;
initial mem[47] = 16'he140;
initial mem[48] = 16'h3041;
initial mem[49] = 16'h1200;
initial mem[50] = 16'he140;
initial mem[51] = 16'h3041;
initial mem[52] = 16'h1200;
initial mem[53] = 16'he141;
initial mem[54] = 16'h3043;
initial mem[55] = 16'h1200;
initial mem[56] = 16'he142;
initial mem[57] = 16'h1004;
initial mem[58] = 16'h4603;
initial mem[59] = 16'h7021;
initial mem[60] = 16'h6f00;
initial mem[61] = 16'h7064;
initial mem[62] = 16'h60f0;
initial mem[63] = 16'h7064;
initial mem[64] = 16'h600f;
initial mem[65] = 16'h7064;
initial mem[66] = 16'h1001;
initial mem[67] = 16'h1006;
initial mem[68] = 16'h3029;
initial mem[69] = 16'hc410;
initial mem[70] = 16'h3121;
initial mem[71] = 16'h2611;
initial mem[72] = 16'h1005;
initial mem[73] = 16'h4003;
initial mem[74] = 16'h1000;
initial mem[75] = 16'he110;
initial mem[76] = 16'h1000;
initial mem[77] = 16'he031;
initial mem[78] = 16'h3d31;
initial mem[79] = 16'h1004;
initial mem[80] = 16'h400c;
initial mem[81] = 16'h1004;
initial mem[82] = 16'h4605;
initial mem[83] = 16'h3011;
initial mem[84] = 16'h1700;
initial mem[85] = 16'he110;
initial mem[86] = 16'h0601;
initial mem[87] = 16'h1fff;
initial mem[88] = 16'h303f;
initial mem[89] = 16'h1002;
initial mem[90] = 16'h3040;
initial mem[91] = 16'h3341;
initial mem[92] = 16'h1005;
initial mem[93] = 16'h410b;
initial mem[94] = 16'h3331;
initial mem[95] = 16'h1005;
initial mem[96] = 16'h4109;
initial mem[97] = 16'h1002;
initial mem[98] = 16'h301e;
initial mem[99] = 16'h1000;
initial mem[100] = 16'he110;
initial mem[101] = 16'h1005;
initial mem[102] = 16'h4607;
initial mem[103] = 16'h1005;
initial mem[104] = 16'h4607;
initial mem[105] = 16'h0048;
initial mem[106] = 16'h0065;
initial mem[107] = 16'h006c;
initial mem[108] = 16'h006c;
initial mem[109] = 16'h006f;
initial mem[110] = 16'h0020;
initial mem[111] = 16'h0077;
initial mem[112] = 16'h006f;
initial mem[113] = 16'h0072;
initial mem[114] = 16'h006c;
initial mem[115] = 16'h0064;
initial mem[116] = 16'h0021;
initial mem[117] = 16'h000d;
initial mem[118] = 16'h000a;
initial mem[119] = 16'h0000;
initial mem[120] = 16'h1002;
initial mem[121] = 16'h3071;
initial mem[122] = 16'h1000;
initial mem[123] = 16'he170;
initial mem[124] = 16'h301f;
initial mem[125] = 16'h1700;
initial mem[126] = 16'he111;
initial mem[127] = 16'h0101;
initial mem[128] = 16'h0000;
initial mem[129] = 16'h0000;
initial mem[130] = 16'h0000;
initial mem[131] = 16'h0000;
initial mem[132] = 16'h0000;
initial mem[133] = 16'h0000;
initial mem[134] = 16'h0000;
initial mem[135] = 16'h0000;
initial mem[136] = 16'h0000;
initial mem[137] = 16'h0000;
initial mem[138] = 16'h0000;
initial mem[139] = 16'h0000;
initial mem[140] = 16'h0000;
initial mem[141] = 16'h0000;
initial mem[142] = 16'h0000;
initial mem[143] = 16'h0000;
initial mem[144] = 16'h0000;
initial mem[145] = 16'h0000;
initial mem[146] = 16'h0000;
initial mem[147] = 16'h0000;
initial mem[148] = 16'h0000;
initial mem[149] = 16'h0000;
initial mem[150] = 16'h0000;
initial mem[151] = 16'h0000;
initial mem[152] = 16'h0000;
initial mem[153] = 16'h0000;
initial mem[154] = 16'h0000;
initial mem[155] = 16'h0000;
initial mem[156] = 16'h0000;
initial mem[157] = 16'h0000;
initial mem[158] = 16'h0000;
initial mem[159] = 16'h0000;
initial mem[160] = 16'h0000;
initial mem[161] = 16'h0000;
initial mem[162] = 16'h0000;
initial mem[163] = 16'h0000;
initial mem[164] = 16'h0000;
initial mem[165] = 16'h0000;
initial mem[166] = 16'h0000;
initial mem[167] = 16'h0000;
initial mem[168] = 16'h0000;
initial mem[169] = 16'h0000;
initial mem[170] = 16'h0000;
initial mem[171] = 16'h0000;
initial mem[172] = 16'h0000;
initial mem[173] = 16'h0000;
initial mem[174] = 16'h0000;
initial mem[175] = 16'h0000;
initial mem[176] = 16'h0000;
initial mem[177] = 16'h0000;
initial mem[178] = 16'h0000;
initial mem[179] = 16'h0000;
initial mem[180] = 16'h0000;
initial mem[181] = 16'h0000;
initial mem[182] = 16'h0000;
initial mem[183] = 16'h0000;
initial mem[184] = 16'h0000;
initial mem[185] = 16'h0000;
initial mem[186] = 16'h0000;
initial mem[187] = 16'h0000;
initial mem[188] = 16'h0000;
initial mem[189] = 16'h0000;
initial mem[190] = 16'h0000;
initial mem[191] = 16'h0000;
initial mem[192] = 16'h0000;
initial mem[193] = 16'h0000;
initial mem[194] = 16'h0000;
initial mem[195] = 16'h0000;
initial mem[196] = 16'h0000;
initial mem[197] = 16'h0000;
initial mem[198] = 16'h0000;
initial mem[199] = 16'h0000;
initial mem[200] = 16'h0000;
initial mem[201] = 16'h0000;
initial mem[202] = 16'h0000;
initial mem[203] = 16'h0000;
initial mem[204] = 16'h0000;
initial mem[205] = 16'h0000;
initial mem[206] = 16'h0000;
initial mem[207] = 16'h0000;
initial mem[208] = 16'h0000;
initial mem[209] = 16'h0000;
initial mem[210] = 16'h0000;
initial mem[211] = 16'h0000;
initial mem[212] = 16'h0000;
initial mem[213] = 16'h0000;
initial mem[214] = 16'h0000;
initial mem[215] = 16'h0000;
initial mem[216] = 16'h0000;
initial mem[217] = 16'h0000;
initial mem[218] = 16'h0000;
initial mem[219] = 16'h0000;
initial mem[220] = 16'h0000;
initial mem[221] = 16'h0000;
initial mem[222] = 16'h0000;
initial mem[223] = 16'h0000;
initial mem[224] = 16'h0000;
initial mem[225] = 16'h0000;
initial mem[226] = 16'h0000;
initial mem[227] = 16'h0000;
initial mem[228] = 16'h0000;
initial mem[229] = 16'h0000;
initial mem[230] = 16'h0000;
initial mem[231] = 16'h0000;
initial mem[232] = 16'h0000;
initial mem[233] = 16'h0000;
initial mem[234] = 16'h0000;
initial mem[235] = 16'h0000;
initial mem[236] = 16'h0000;
initial mem[237] = 16'h0000;
initial mem[238] = 16'h0000;
initial mem[239] = 16'h0000;
initial mem[240] = 16'h0000;
initial mem[241] = 16'h0000;
initial mem[242] = 16'h0000;
initial mem[243] = 16'h0000;
initial mem[244] = 16'h0000;
initial mem[245] = 16'h0000;
initial mem[246] = 16'h0000;
initial mem[247] = 16'h0000;
initial mem[248] = 16'h0000;
initial mem[249] = 16'h0000;
initial mem[250] = 16'h0000;
initial mem[251] = 16'h0000;
initial mem[252] = 16'h0000;
initial mem[253] = 16'h0000;
initial mem[254] = 16'h0000;
initial mem[255] = 16'h0000;
always @(posedge CLK)
begin
       dout <= mem[ADDRESS];
end
endmodule
