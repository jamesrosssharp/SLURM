/* rom.v : rom */

module rom
#(parameter BITS = 16, ADDRESS_BITS = 16)
(
	input CLK,
	input [ADDRESS_BITS - 1 : 0]  ADDRESS,
	output [BITS - 1 : 0] DATA_OUT,
);

localparam ROM_ADDRESS_BITS = 12;

reg [BITS - 1:0] mem [(1 << ROM_ADDRESS_BITS) - 1:0];
reg [BITS - 1:0] dout;
assign DATA_OUT = dout;
initial mem[0] = 16'h0000;
initial mem[1] = 16'h1fff;
initial mem[2] = 16'h306f;
initial mem[3] = 16'h3002;
initial mem[4] = 16'h1140;
initial mem[5] = 16'h6102;
initial mem[6] = 16'h1001;
initial mem[7] = 16'h3044;
initial mem[8] = 16'h1fff;
initial mem[9] = 16'h303f;
initial mem[10] = 16'h3331;
initial mem[11] = 16'h1000;
initial mem[12] = 16'h410a;
initial mem[13] = 16'h3341;
initial mem[14] = 16'h1000;
initial mem[15] = 16'h4108;
initial mem[16] = 16'h1400;
initial mem[17] = 16'h30b0;
initial mem[18] = 16'h3161;
initial mem[19] = 16'h2006;
initial mem[20] = 16'h3018;
initial mem[21] = 16'h1140;
initial mem[22] = 16'h6100;
initial mem[23] = 16'h1140;
initial mem[24] = 16'h6111;
initial mem[25] = 16'h3001;
initial mem[26] = 16'h1140;
initial mem[27] = 16'h6102;
initial mem[28] = 16'h1140;
initial mem[29] = 16'h6004;
initial mem[30] = 16'h3d01;
initial mem[31] = 16'h1001;
initial mem[32] = 16'h400c;
initial mem[33] = 16'h1140;
initial mem[34] = 16'h6003;
initial mem[35] = 16'h570b;
initial mem[36] = 16'h020b;
initial mem[37] = 16'h26bb;
initial mem[38] = 16'h1400;
initial mem[39] = 16'h4000;
initial mem[40] = 16'h1001;
initial mem[41] = 16'h4602;
initial mem[42] = 16'h0000;
initial mem[43] = 16'h0000;
initial mem[44] = 16'h0000;
initial mem[45] = 16'h0000;
initial mem[46] = 16'h0000;
initial mem[47] = 16'h0000;
initial mem[48] = 16'h0000;
initial mem[49] = 16'h0000;
initial mem[50] = 16'h0000;
initial mem[51] = 16'h0000;
initial mem[52] = 16'h0000;
initial mem[53] = 16'h0000;
initial mem[54] = 16'h0000;
initial mem[55] = 16'h0000;
initial mem[56] = 16'h0000;
initial mem[57] = 16'h0000;
initial mem[58] = 16'h0000;
initial mem[59] = 16'h0000;
initial mem[60] = 16'h0000;
initial mem[61] = 16'h0000;
initial mem[62] = 16'h0000;
initial mem[63] = 16'h0000;
initial mem[64] = 16'h0000;
initial mem[65] = 16'h0000;
initial mem[66] = 16'h0000;
initial mem[67] = 16'h0000;
initial mem[68] = 16'h0000;
initial mem[69] = 16'h0000;
initial mem[70] = 16'h0000;
initial mem[71] = 16'h0000;
initial mem[72] = 16'h0000;
initial mem[73] = 16'h0000;
initial mem[74] = 16'h0000;
initial mem[75] = 16'h0000;
initial mem[76] = 16'h0000;
initial mem[77] = 16'h0000;
initial mem[78] = 16'h0000;
initial mem[79] = 16'h0000;
initial mem[80] = 16'h0000;
initial mem[81] = 16'h0000;
initial mem[82] = 16'h0000;
initial mem[83] = 16'h0000;
initial mem[84] = 16'h0000;
initial mem[85] = 16'h0000;
initial mem[86] = 16'h0000;
initial mem[87] = 16'h0000;
initial mem[88] = 16'h0000;
initial mem[89] = 16'h0000;
initial mem[90] = 16'h0000;
initial mem[91] = 16'h0000;
initial mem[92] = 16'h0000;
initial mem[93] = 16'h0000;
initial mem[94] = 16'h0000;
initial mem[95] = 16'h0000;
initial mem[96] = 16'h0000;
initial mem[97] = 16'h0000;
initial mem[98] = 16'h0000;
initial mem[99] = 16'h0000;
initial mem[100] = 16'h0000;
initial mem[101] = 16'h0000;
initial mem[102] = 16'h0000;
initial mem[103] = 16'h0000;
initial mem[104] = 16'h0000;
initial mem[105] = 16'h0000;
initial mem[106] = 16'h0000;
initial mem[107] = 16'h0000;
initial mem[108] = 16'h0000;
initial mem[109] = 16'h0000;
initial mem[110] = 16'h0000;
initial mem[111] = 16'h0000;
initial mem[112] = 16'h0000;
initial mem[113] = 16'h0000;
initial mem[114] = 16'h0000;
initial mem[115] = 16'h0000;
initial mem[116] = 16'h0000;
initial mem[117] = 16'h0000;
initial mem[118] = 16'h0000;
initial mem[119] = 16'h0000;
initial mem[120] = 16'h0000;
initial mem[121] = 16'h0000;
initial mem[122] = 16'h0000;
initial mem[123] = 16'h0000;
initial mem[124] = 16'h0000;
initial mem[125] = 16'h0000;
initial mem[126] = 16'h0000;
initial mem[127] = 16'h0000;
initial mem[128] = 16'h0000;
initial mem[129] = 16'h0000;
initial mem[130] = 16'h0000;
initial mem[131] = 16'h0000;
initial mem[132] = 16'h0000;
initial mem[133] = 16'h0000;
initial mem[134] = 16'h0000;
initial mem[135] = 16'h0000;
initial mem[136] = 16'h0000;
initial mem[137] = 16'h0000;
initial mem[138] = 16'h0000;
initial mem[139] = 16'h0000;
initial mem[140] = 16'h0000;
initial mem[141] = 16'h0000;
initial mem[142] = 16'h0000;
initial mem[143] = 16'h0000;
initial mem[144] = 16'h0000;
initial mem[145] = 16'h0000;
initial mem[146] = 16'h0000;
initial mem[147] = 16'h0000;
initial mem[148] = 16'h0000;
initial mem[149] = 16'h0000;
initial mem[150] = 16'h0000;
initial mem[151] = 16'h0000;
initial mem[152] = 16'h0000;
initial mem[153] = 16'h0000;
initial mem[154] = 16'h0000;
initial mem[155] = 16'h0000;
initial mem[156] = 16'h0000;
initial mem[157] = 16'h0000;
initial mem[158] = 16'h0000;
initial mem[159] = 16'h0000;
initial mem[160] = 16'h0000;
initial mem[161] = 16'h0000;
initial mem[162] = 16'h0000;
initial mem[163] = 16'h0000;
initial mem[164] = 16'h0000;
initial mem[165] = 16'h0000;
initial mem[166] = 16'h0000;
initial mem[167] = 16'h0000;
initial mem[168] = 16'h0000;
initial mem[169] = 16'h0000;
initial mem[170] = 16'h0000;
initial mem[171] = 16'h0000;
initial mem[172] = 16'h0000;
initial mem[173] = 16'h0000;
initial mem[174] = 16'h0000;
initial mem[175] = 16'h0000;
initial mem[176] = 16'h0000;
initial mem[177] = 16'h0000;
initial mem[178] = 16'h0000;
initial mem[179] = 16'h0000;
initial mem[180] = 16'h0000;
initial mem[181] = 16'h0000;
initial mem[182] = 16'h0000;
initial mem[183] = 16'h0000;
initial mem[184] = 16'h0000;
initial mem[185] = 16'h0000;
initial mem[186] = 16'h0000;
initial mem[187] = 16'h0000;
initial mem[188] = 16'h0000;
initial mem[189] = 16'h0000;
initial mem[190] = 16'h0000;
initial mem[191] = 16'h0000;
initial mem[192] = 16'h0000;
initial mem[193] = 16'h0000;
initial mem[194] = 16'h0000;
initial mem[195] = 16'h0000;
initial mem[196] = 16'h0000;
initial mem[197] = 16'h0000;
initial mem[198] = 16'h0000;
initial mem[199] = 16'h0000;
initial mem[200] = 16'h0000;
initial mem[201] = 16'h0000;
initial mem[202] = 16'h0000;
initial mem[203] = 16'h0000;
initial mem[204] = 16'h0000;
initial mem[205] = 16'h0000;
initial mem[206] = 16'h0000;
initial mem[207] = 16'h0000;
initial mem[208] = 16'h0000;
initial mem[209] = 16'h0000;
initial mem[210] = 16'h0000;
initial mem[211] = 16'h0000;
initial mem[212] = 16'h0000;
initial mem[213] = 16'h0000;
initial mem[214] = 16'h0000;
initial mem[215] = 16'h0000;
initial mem[216] = 16'h0000;
initial mem[217] = 16'h0000;
initial mem[218] = 16'h0000;
initial mem[219] = 16'h0000;
initial mem[220] = 16'h0000;
initial mem[221] = 16'h0000;
initial mem[222] = 16'h0000;
initial mem[223] = 16'h0000;
initial mem[224] = 16'h0000;
initial mem[225] = 16'h0000;
initial mem[226] = 16'h0000;
initial mem[227] = 16'h0000;
initial mem[228] = 16'h0000;
initial mem[229] = 16'h0000;
initial mem[230] = 16'h0000;
initial mem[231] = 16'h0000;
initial mem[232] = 16'h0000;
initial mem[233] = 16'h0000;
initial mem[234] = 16'h0000;
initial mem[235] = 16'h0000;
initial mem[236] = 16'h0000;
initial mem[237] = 16'h0000;
initial mem[238] = 16'h0000;
initial mem[239] = 16'h0000;
initial mem[240] = 16'h0000;
initial mem[241] = 16'h0000;
initial mem[242] = 16'h0000;
initial mem[243] = 16'h0000;
initial mem[244] = 16'h0000;
initial mem[245] = 16'h0000;
initial mem[246] = 16'h0000;
initial mem[247] = 16'h0000;
initial mem[248] = 16'h0000;
initial mem[249] = 16'h0000;
initial mem[250] = 16'h0000;
initial mem[251] = 16'h0000;
initial mem[252] = 16'h0000;
initial mem[253] = 16'h0000;
initial mem[254] = 16'h0000;
initial mem[255] = 16'h0000;
initial mem[256] = 16'h0000;
initial mem[257] = 16'h0000;
initial mem[258] = 16'h0000;
initial mem[259] = 16'h0000;
initial mem[260] = 16'h0000;
initial mem[261] = 16'h0000;
initial mem[262] = 16'h0000;
initial mem[263] = 16'h0000;
initial mem[264] = 16'h0000;
initial mem[265] = 16'h0000;
initial mem[266] = 16'h0000;
initial mem[267] = 16'h0000;
initial mem[268] = 16'h0000;
initial mem[269] = 16'h0000;
initial mem[270] = 16'h0000;
initial mem[271] = 16'h0000;
initial mem[272] = 16'h0000;
initial mem[273] = 16'h0000;
initial mem[274] = 16'h0000;
initial mem[275] = 16'h0000;
initial mem[276] = 16'h0000;
initial mem[277] = 16'h0000;
initial mem[278] = 16'h0000;
initial mem[279] = 16'h0000;
initial mem[280] = 16'h0000;
initial mem[281] = 16'h0000;
initial mem[282] = 16'h0000;
initial mem[283] = 16'h0000;
initial mem[284] = 16'h0000;
initial mem[285] = 16'h0000;
initial mem[286] = 16'h0000;
initial mem[287] = 16'h0000;
initial mem[288] = 16'h0000;
initial mem[289] = 16'h0000;
initial mem[290] = 16'h0000;
initial mem[291] = 16'h0000;
initial mem[292] = 16'h0000;
initial mem[293] = 16'h0000;
initial mem[294] = 16'h0000;
initial mem[295] = 16'h0000;
initial mem[296] = 16'h0000;
initial mem[297] = 16'h0000;
initial mem[298] = 16'h0000;
initial mem[299] = 16'h0000;
initial mem[300] = 16'h0000;
initial mem[301] = 16'h0000;
initial mem[302] = 16'h0000;
initial mem[303] = 16'h0000;
initial mem[304] = 16'h0000;
initial mem[305] = 16'h0000;
initial mem[306] = 16'h0000;
initial mem[307] = 16'h0000;
initial mem[308] = 16'h0000;
initial mem[309] = 16'h0000;
initial mem[310] = 16'h0000;
initial mem[311] = 16'h0000;
initial mem[312] = 16'h0000;
initial mem[313] = 16'h0000;
initial mem[314] = 16'h0000;
initial mem[315] = 16'h0000;
initial mem[316] = 16'h0000;
initial mem[317] = 16'h0000;
initial mem[318] = 16'h0000;
initial mem[319] = 16'h0000;
initial mem[320] = 16'h0000;
initial mem[321] = 16'h0000;
initial mem[322] = 16'h0000;
initial mem[323] = 16'h0000;
initial mem[324] = 16'h0000;
initial mem[325] = 16'h0000;
initial mem[326] = 16'h0000;
initial mem[327] = 16'h0000;
initial mem[328] = 16'h0000;
initial mem[329] = 16'h0000;
initial mem[330] = 16'h0000;
initial mem[331] = 16'h0000;
initial mem[332] = 16'h0000;
initial mem[333] = 16'h0000;
initial mem[334] = 16'h0000;
initial mem[335] = 16'h0000;
initial mem[336] = 16'h0000;
initial mem[337] = 16'h0000;
initial mem[338] = 16'h0000;
initial mem[339] = 16'h0000;
initial mem[340] = 16'h0000;
initial mem[341] = 16'h0000;
initial mem[342] = 16'h0000;
initial mem[343] = 16'h0000;
initial mem[344] = 16'h0000;
initial mem[345] = 16'h0000;
initial mem[346] = 16'h0000;
initial mem[347] = 16'h0000;
initial mem[348] = 16'h0000;
initial mem[349] = 16'h0000;
initial mem[350] = 16'h0000;
initial mem[351] = 16'h0000;
initial mem[352] = 16'h0000;
initial mem[353] = 16'h0000;
initial mem[354] = 16'h0000;
initial mem[355] = 16'h0000;
initial mem[356] = 16'h0000;
initial mem[357] = 16'h0000;
initial mem[358] = 16'h0000;
initial mem[359] = 16'h0000;
initial mem[360] = 16'h0000;
initial mem[361] = 16'h0000;
initial mem[362] = 16'h0000;
initial mem[363] = 16'h0000;
initial mem[364] = 16'h0000;
initial mem[365] = 16'h0000;
initial mem[366] = 16'h0000;
initial mem[367] = 16'h0000;
initial mem[368] = 16'h0000;
initial mem[369] = 16'h0000;
initial mem[370] = 16'h0000;
initial mem[371] = 16'h0000;
initial mem[372] = 16'h0000;
initial mem[373] = 16'h0000;
initial mem[374] = 16'h0000;
initial mem[375] = 16'h0000;
initial mem[376] = 16'h0000;
initial mem[377] = 16'h0000;
initial mem[378] = 16'h0000;
initial mem[379] = 16'h0000;
initial mem[380] = 16'h0000;
initial mem[381] = 16'h0000;
initial mem[382] = 16'h0000;
initial mem[383] = 16'h0000;
initial mem[384] = 16'h0000;
initial mem[385] = 16'h0000;
initial mem[386] = 16'h0000;
initial mem[387] = 16'h0000;
initial mem[388] = 16'h0000;
initial mem[389] = 16'h0000;
initial mem[390] = 16'h0000;
initial mem[391] = 16'h0000;
initial mem[392] = 16'h0000;
initial mem[393] = 16'h0000;
initial mem[394] = 16'h0000;
initial mem[395] = 16'h0000;
initial mem[396] = 16'h0000;
initial mem[397] = 16'h0000;
initial mem[398] = 16'h0000;
initial mem[399] = 16'h0000;
initial mem[400] = 16'h0000;
initial mem[401] = 16'h0000;
initial mem[402] = 16'h0000;
initial mem[403] = 16'h0000;
initial mem[404] = 16'h0000;
initial mem[405] = 16'h0000;
initial mem[406] = 16'h0000;
initial mem[407] = 16'h0000;
initial mem[408] = 16'h0000;
initial mem[409] = 16'h0000;
initial mem[410] = 16'h0000;
initial mem[411] = 16'h0000;
initial mem[412] = 16'h0000;
initial mem[413] = 16'h0000;
initial mem[414] = 16'h0000;
initial mem[415] = 16'h0000;
initial mem[416] = 16'h0000;
initial mem[417] = 16'h0000;
initial mem[418] = 16'h0000;
initial mem[419] = 16'h0000;
initial mem[420] = 16'h0000;
initial mem[421] = 16'h0000;
initial mem[422] = 16'h0000;
initial mem[423] = 16'h0000;
initial mem[424] = 16'h0000;
initial mem[425] = 16'h0000;
initial mem[426] = 16'h0000;
initial mem[427] = 16'h0000;
initial mem[428] = 16'h0000;
initial mem[429] = 16'h0000;
initial mem[430] = 16'h0000;
initial mem[431] = 16'h0000;
initial mem[432] = 16'h0000;
initial mem[433] = 16'h0000;
initial mem[434] = 16'h0000;
initial mem[435] = 16'h0000;
initial mem[436] = 16'h0000;
initial mem[437] = 16'h0000;
initial mem[438] = 16'h0000;
initial mem[439] = 16'h0000;
initial mem[440] = 16'h0000;
initial mem[441] = 16'h0000;
initial mem[442] = 16'h0000;
initial mem[443] = 16'h0000;
initial mem[444] = 16'h0000;
initial mem[445] = 16'h0000;
initial mem[446] = 16'h0000;
initial mem[447] = 16'h0000;
initial mem[448] = 16'h0000;
initial mem[449] = 16'h0000;
initial mem[450] = 16'h0000;
initial mem[451] = 16'h0000;
initial mem[452] = 16'h0000;
initial mem[453] = 16'h0000;
initial mem[454] = 16'h0000;
initial mem[455] = 16'h0000;
initial mem[456] = 16'h0000;
initial mem[457] = 16'h0000;
initial mem[458] = 16'h0000;
initial mem[459] = 16'h0000;
initial mem[460] = 16'h0000;
initial mem[461] = 16'h0000;
initial mem[462] = 16'h0000;
initial mem[463] = 16'h0000;
initial mem[464] = 16'h0000;
initial mem[465] = 16'h0000;
initial mem[466] = 16'h0000;
initial mem[467] = 16'h0000;
initial mem[468] = 16'h0000;
initial mem[469] = 16'h0000;
initial mem[470] = 16'h0000;
initial mem[471] = 16'h0000;
initial mem[472] = 16'h0000;
initial mem[473] = 16'h0000;
initial mem[474] = 16'h0000;
initial mem[475] = 16'h0000;
initial mem[476] = 16'h0000;
initial mem[477] = 16'h0000;
initial mem[478] = 16'h0000;
initial mem[479] = 16'h0000;
initial mem[480] = 16'h0000;
initial mem[481] = 16'h0000;
initial mem[482] = 16'h0000;
initial mem[483] = 16'h0000;
initial mem[484] = 16'h0000;
initial mem[485] = 16'h0000;
initial mem[486] = 16'h0000;
initial mem[487] = 16'h0000;
initial mem[488] = 16'h0000;
initial mem[489] = 16'h0000;
initial mem[490] = 16'h0000;
initial mem[491] = 16'h0000;
initial mem[492] = 16'h0000;
initial mem[493] = 16'h0000;
initial mem[494] = 16'h0000;
initial mem[495] = 16'h0000;
initial mem[496] = 16'h0000;
initial mem[497] = 16'h0000;
initial mem[498] = 16'h0000;
initial mem[499] = 16'h0000;
initial mem[500] = 16'h0000;
initial mem[501] = 16'h0000;
initial mem[502] = 16'h0000;
initial mem[503] = 16'h0000;
initial mem[504] = 16'h0000;
initial mem[505] = 16'h0000;
initial mem[506] = 16'h0000;
initial mem[507] = 16'h0000;
initial mem[508] = 16'h0000;
initial mem[509] = 16'h0000;
initial mem[510] = 16'h0000;
initial mem[511] = 16'h0000;
initial mem[512] = 16'h0000;
initial mem[513] = 16'h0000;
initial mem[514] = 16'h0000;
initial mem[515] = 16'h0000;
initial mem[516] = 16'h0000;
initial mem[517] = 16'h0000;
initial mem[518] = 16'h0000;
initial mem[519] = 16'h0000;
initial mem[520] = 16'h0000;
initial mem[521] = 16'h0000;
initial mem[522] = 16'h0000;
initial mem[523] = 16'h0000;
initial mem[524] = 16'h0000;
initial mem[525] = 16'h0000;
initial mem[526] = 16'h0000;
initial mem[527] = 16'h0000;
initial mem[528] = 16'h0000;
initial mem[529] = 16'h0000;
initial mem[530] = 16'h0000;
initial mem[531] = 16'h0000;
initial mem[532] = 16'h0000;
initial mem[533] = 16'h0000;
initial mem[534] = 16'h0000;
initial mem[535] = 16'h0000;
initial mem[536] = 16'h0000;
initial mem[537] = 16'h0000;
initial mem[538] = 16'h0000;
initial mem[539] = 16'h0000;
initial mem[540] = 16'h0000;
initial mem[541] = 16'h0000;
initial mem[542] = 16'h0000;
initial mem[543] = 16'h0000;
initial mem[544] = 16'h0000;
initial mem[545] = 16'h0000;
initial mem[546] = 16'h0000;
initial mem[547] = 16'h0000;
initial mem[548] = 16'h0000;
initial mem[549] = 16'h0000;
initial mem[550] = 16'h0000;
initial mem[551] = 16'h0000;
initial mem[552] = 16'h0000;
initial mem[553] = 16'h0000;
initial mem[554] = 16'h0000;
initial mem[555] = 16'h0000;
initial mem[556] = 16'h0000;
initial mem[557] = 16'h0000;
initial mem[558] = 16'h0000;
initial mem[559] = 16'h0000;
initial mem[560] = 16'h0000;
initial mem[561] = 16'h0000;
initial mem[562] = 16'h0000;
initial mem[563] = 16'h0000;
initial mem[564] = 16'h0000;
initial mem[565] = 16'h0000;
initial mem[566] = 16'h0000;
initial mem[567] = 16'h0000;
initial mem[568] = 16'h0000;
initial mem[569] = 16'h0000;
initial mem[570] = 16'h0000;
initial mem[571] = 16'h0000;
initial mem[572] = 16'h0000;
initial mem[573] = 16'h0000;
initial mem[574] = 16'h0000;
initial mem[575] = 16'h0000;
initial mem[576] = 16'h0000;
initial mem[577] = 16'h0000;
initial mem[578] = 16'h0000;
initial mem[579] = 16'h0000;
initial mem[580] = 16'h0000;
initial mem[581] = 16'h0000;
initial mem[582] = 16'h0000;
initial mem[583] = 16'h0000;
initial mem[584] = 16'h0000;
initial mem[585] = 16'h0000;
initial mem[586] = 16'h0000;
initial mem[587] = 16'h0000;
initial mem[588] = 16'h0000;
initial mem[589] = 16'h0000;
initial mem[590] = 16'h0000;
initial mem[591] = 16'h0000;
initial mem[592] = 16'h0000;
initial mem[593] = 16'h0000;
initial mem[594] = 16'h0000;
initial mem[595] = 16'h0000;
initial mem[596] = 16'h0000;
initial mem[597] = 16'h0000;
initial mem[598] = 16'h0000;
initial mem[599] = 16'h0000;
initial mem[600] = 16'h0000;
initial mem[601] = 16'h0000;
initial mem[602] = 16'h0000;
initial mem[603] = 16'h0000;
initial mem[604] = 16'h0000;
initial mem[605] = 16'h0000;
initial mem[606] = 16'h0000;
initial mem[607] = 16'h0000;
initial mem[608] = 16'h0000;
initial mem[609] = 16'h0000;
initial mem[610] = 16'h0000;
initial mem[611] = 16'h0000;
initial mem[612] = 16'h0000;
initial mem[613] = 16'h0000;
initial mem[614] = 16'h0000;
initial mem[615] = 16'h0000;
initial mem[616] = 16'h0000;
initial mem[617] = 16'h0000;
initial mem[618] = 16'h0000;
initial mem[619] = 16'h0000;
initial mem[620] = 16'h0000;
initial mem[621] = 16'h0000;
initial mem[622] = 16'h0000;
initial mem[623] = 16'h0000;
initial mem[624] = 16'h0000;
initial mem[625] = 16'h0000;
initial mem[626] = 16'h0000;
initial mem[627] = 16'h0000;
initial mem[628] = 16'h0000;
initial mem[629] = 16'h0000;
initial mem[630] = 16'h0000;
initial mem[631] = 16'h0000;
initial mem[632] = 16'h0000;
initial mem[633] = 16'h0000;
initial mem[634] = 16'h0000;
initial mem[635] = 16'h0000;
initial mem[636] = 16'h0000;
initial mem[637] = 16'h0000;
initial mem[638] = 16'h0000;
initial mem[639] = 16'h0000;
initial mem[640] = 16'h0000;
initial mem[641] = 16'h0000;
initial mem[642] = 16'h0000;
initial mem[643] = 16'h0000;
initial mem[644] = 16'h0000;
initial mem[645] = 16'h0000;
initial mem[646] = 16'h0000;
initial mem[647] = 16'h0000;
initial mem[648] = 16'h0000;
initial mem[649] = 16'h0000;
initial mem[650] = 16'h0000;
initial mem[651] = 16'h0000;
initial mem[652] = 16'h0000;
initial mem[653] = 16'h0000;
initial mem[654] = 16'h0000;
initial mem[655] = 16'h0000;
initial mem[656] = 16'h0000;
initial mem[657] = 16'h0000;
initial mem[658] = 16'h0000;
initial mem[659] = 16'h0000;
initial mem[660] = 16'h0000;
initial mem[661] = 16'h0000;
initial mem[662] = 16'h0000;
initial mem[663] = 16'h0000;
initial mem[664] = 16'h0000;
initial mem[665] = 16'h0000;
initial mem[666] = 16'h0000;
initial mem[667] = 16'h0000;
initial mem[668] = 16'h0000;
initial mem[669] = 16'h0000;
initial mem[670] = 16'h0000;
initial mem[671] = 16'h0000;
initial mem[672] = 16'h0000;
initial mem[673] = 16'h0000;
initial mem[674] = 16'h0000;
initial mem[675] = 16'h0000;
initial mem[676] = 16'h0000;
initial mem[677] = 16'h0000;
initial mem[678] = 16'h0000;
initial mem[679] = 16'h0000;
initial mem[680] = 16'h0000;
initial mem[681] = 16'h0000;
initial mem[682] = 16'h0000;
initial mem[683] = 16'h0000;
initial mem[684] = 16'h0000;
initial mem[685] = 16'h0000;
initial mem[686] = 16'h0000;
initial mem[687] = 16'h0000;
initial mem[688] = 16'h0000;
initial mem[689] = 16'h0000;
initial mem[690] = 16'h0000;
initial mem[691] = 16'h0000;
initial mem[692] = 16'h0000;
initial mem[693] = 16'h0000;
initial mem[694] = 16'h0000;
initial mem[695] = 16'h0000;
initial mem[696] = 16'h0000;
initial mem[697] = 16'h0000;
initial mem[698] = 16'h0000;
initial mem[699] = 16'h0000;
initial mem[700] = 16'h0000;
initial mem[701] = 16'h0000;
initial mem[702] = 16'h0000;
initial mem[703] = 16'h0000;
initial mem[704] = 16'h0000;
initial mem[705] = 16'h0000;
initial mem[706] = 16'h0000;
initial mem[707] = 16'h0000;
initial mem[708] = 16'h0000;
initial mem[709] = 16'h0000;
initial mem[710] = 16'h0000;
initial mem[711] = 16'h0000;
initial mem[712] = 16'h0000;
initial mem[713] = 16'h0000;
initial mem[714] = 16'h0000;
initial mem[715] = 16'h0000;
initial mem[716] = 16'h0000;
initial mem[717] = 16'h0000;
initial mem[718] = 16'h0000;
initial mem[719] = 16'h0000;
initial mem[720] = 16'h0000;
initial mem[721] = 16'h0000;
initial mem[722] = 16'h0000;
initial mem[723] = 16'h0000;
initial mem[724] = 16'h0000;
initial mem[725] = 16'h0000;
initial mem[726] = 16'h0000;
initial mem[727] = 16'h0000;
initial mem[728] = 16'h0000;
initial mem[729] = 16'h0000;
initial mem[730] = 16'h0000;
initial mem[731] = 16'h0000;
initial mem[732] = 16'h0000;
initial mem[733] = 16'h0000;
initial mem[734] = 16'h0000;
initial mem[735] = 16'h0000;
initial mem[736] = 16'h0000;
initial mem[737] = 16'h0000;
initial mem[738] = 16'h0000;
initial mem[739] = 16'h0000;
initial mem[740] = 16'h0000;
initial mem[741] = 16'h0000;
initial mem[742] = 16'h0000;
initial mem[743] = 16'h0000;
initial mem[744] = 16'h0000;
initial mem[745] = 16'h0000;
initial mem[746] = 16'h0000;
initial mem[747] = 16'h0000;
initial mem[748] = 16'h0000;
initial mem[749] = 16'h0000;
initial mem[750] = 16'h0000;
initial mem[751] = 16'h0000;
initial mem[752] = 16'h0000;
initial mem[753] = 16'h0000;
initial mem[754] = 16'h0000;
initial mem[755] = 16'h0000;
initial mem[756] = 16'h0000;
initial mem[757] = 16'h0000;
initial mem[758] = 16'h0000;
initial mem[759] = 16'h0000;
initial mem[760] = 16'h0000;
initial mem[761] = 16'h0000;
initial mem[762] = 16'h0000;
initial mem[763] = 16'h0000;
initial mem[764] = 16'h0000;
initial mem[765] = 16'h0000;
initial mem[766] = 16'h0000;
initial mem[767] = 16'h0000;
initial mem[768] = 16'h0000;
initial mem[769] = 16'h0000;
initial mem[770] = 16'h0000;
initial mem[771] = 16'h0000;
initial mem[772] = 16'h0000;
initial mem[773] = 16'h0000;
initial mem[774] = 16'h0000;
initial mem[775] = 16'h0000;
initial mem[776] = 16'h0000;
initial mem[777] = 16'h0000;
initial mem[778] = 16'h0000;
initial mem[779] = 16'h0000;
initial mem[780] = 16'h0000;
initial mem[781] = 16'h0000;
initial mem[782] = 16'h0000;
initial mem[783] = 16'h0000;
initial mem[784] = 16'h0000;
initial mem[785] = 16'h0000;
initial mem[786] = 16'h0000;
initial mem[787] = 16'h0000;
initial mem[788] = 16'h0000;
initial mem[789] = 16'h0000;
initial mem[790] = 16'h0000;
initial mem[791] = 16'h0000;
initial mem[792] = 16'h0000;
initial mem[793] = 16'h0000;
initial mem[794] = 16'h0000;
initial mem[795] = 16'h0000;
initial mem[796] = 16'h0000;
initial mem[797] = 16'h0000;
initial mem[798] = 16'h0000;
initial mem[799] = 16'h0000;
initial mem[800] = 16'h0000;
initial mem[801] = 16'h0000;
initial mem[802] = 16'h0000;
initial mem[803] = 16'h0000;
initial mem[804] = 16'h0000;
initial mem[805] = 16'h0000;
initial mem[806] = 16'h0000;
initial mem[807] = 16'h0000;
initial mem[808] = 16'h0000;
initial mem[809] = 16'h0000;
initial mem[810] = 16'h0000;
initial mem[811] = 16'h0000;
initial mem[812] = 16'h0000;
initial mem[813] = 16'h0000;
initial mem[814] = 16'h0000;
initial mem[815] = 16'h0000;
initial mem[816] = 16'h0000;
initial mem[817] = 16'h0000;
initial mem[818] = 16'h0000;
initial mem[819] = 16'h0000;
initial mem[820] = 16'h0000;
initial mem[821] = 16'h0000;
initial mem[822] = 16'h0000;
initial mem[823] = 16'h0000;
initial mem[824] = 16'h0000;
initial mem[825] = 16'h0000;
initial mem[826] = 16'h0000;
initial mem[827] = 16'h0000;
initial mem[828] = 16'h0000;
initial mem[829] = 16'h0000;
initial mem[830] = 16'h0000;
initial mem[831] = 16'h0000;
initial mem[832] = 16'h0000;
initial mem[833] = 16'h0000;
initial mem[834] = 16'h0000;
initial mem[835] = 16'h0000;
initial mem[836] = 16'h0000;
initial mem[837] = 16'h0000;
initial mem[838] = 16'h0000;
initial mem[839] = 16'h0000;
initial mem[840] = 16'h0000;
initial mem[841] = 16'h0000;
initial mem[842] = 16'h0000;
initial mem[843] = 16'h0000;
initial mem[844] = 16'h0000;
initial mem[845] = 16'h0000;
initial mem[846] = 16'h0000;
initial mem[847] = 16'h0000;
initial mem[848] = 16'h0000;
initial mem[849] = 16'h0000;
initial mem[850] = 16'h0000;
initial mem[851] = 16'h0000;
initial mem[852] = 16'h0000;
initial mem[853] = 16'h0000;
initial mem[854] = 16'h0000;
initial mem[855] = 16'h0000;
initial mem[856] = 16'h0000;
initial mem[857] = 16'h0000;
initial mem[858] = 16'h0000;
initial mem[859] = 16'h0000;
initial mem[860] = 16'h0000;
initial mem[861] = 16'h0000;
initial mem[862] = 16'h0000;
initial mem[863] = 16'h0000;
initial mem[864] = 16'h0000;
initial mem[865] = 16'h0000;
initial mem[866] = 16'h0000;
initial mem[867] = 16'h0000;
initial mem[868] = 16'h0000;
initial mem[869] = 16'h0000;
initial mem[870] = 16'h0000;
initial mem[871] = 16'h0000;
initial mem[872] = 16'h0000;
initial mem[873] = 16'h0000;
initial mem[874] = 16'h0000;
initial mem[875] = 16'h0000;
initial mem[876] = 16'h0000;
initial mem[877] = 16'h0000;
initial mem[878] = 16'h0000;
initial mem[879] = 16'h0000;
initial mem[880] = 16'h0000;
initial mem[881] = 16'h0000;
initial mem[882] = 16'h0000;
initial mem[883] = 16'h0000;
initial mem[884] = 16'h0000;
initial mem[885] = 16'h0000;
initial mem[886] = 16'h0000;
initial mem[887] = 16'h0000;
initial mem[888] = 16'h0000;
initial mem[889] = 16'h0000;
initial mem[890] = 16'h0000;
initial mem[891] = 16'h0000;
initial mem[892] = 16'h0000;
initial mem[893] = 16'h0000;
initial mem[894] = 16'h0000;
initial mem[895] = 16'h0000;
initial mem[896] = 16'h0000;
initial mem[897] = 16'h0000;
initial mem[898] = 16'h0000;
initial mem[899] = 16'h0000;
initial mem[900] = 16'h0000;
initial mem[901] = 16'h0000;
initial mem[902] = 16'h0000;
initial mem[903] = 16'h0000;
initial mem[904] = 16'h0000;
initial mem[905] = 16'h0000;
initial mem[906] = 16'h0000;
initial mem[907] = 16'h0000;
initial mem[908] = 16'h0000;
initial mem[909] = 16'h0000;
initial mem[910] = 16'h0000;
initial mem[911] = 16'h0000;
initial mem[912] = 16'h0000;
initial mem[913] = 16'h0000;
initial mem[914] = 16'h0000;
initial mem[915] = 16'h0000;
initial mem[916] = 16'h0000;
initial mem[917] = 16'h0000;
initial mem[918] = 16'h0000;
initial mem[919] = 16'h0000;
initial mem[920] = 16'h0000;
initial mem[921] = 16'h0000;
initial mem[922] = 16'h0000;
initial mem[923] = 16'h0000;
initial mem[924] = 16'h0000;
initial mem[925] = 16'h0000;
initial mem[926] = 16'h0000;
initial mem[927] = 16'h0000;
initial mem[928] = 16'h0000;
initial mem[929] = 16'h0000;
initial mem[930] = 16'h0000;
initial mem[931] = 16'h0000;
initial mem[932] = 16'h0000;
initial mem[933] = 16'h0000;
initial mem[934] = 16'h0000;
initial mem[935] = 16'h0000;
initial mem[936] = 16'h0000;
initial mem[937] = 16'h0000;
initial mem[938] = 16'h0000;
initial mem[939] = 16'h0000;
initial mem[940] = 16'h0000;
initial mem[941] = 16'h0000;
initial mem[942] = 16'h0000;
initial mem[943] = 16'h0000;
initial mem[944] = 16'h0000;
initial mem[945] = 16'h0000;
initial mem[946] = 16'h0000;
initial mem[947] = 16'h0000;
initial mem[948] = 16'h0000;
initial mem[949] = 16'h0000;
initial mem[950] = 16'h0000;
initial mem[951] = 16'h0000;
initial mem[952] = 16'h0000;
initial mem[953] = 16'h0000;
initial mem[954] = 16'h0000;
initial mem[955] = 16'h0000;
initial mem[956] = 16'h0000;
initial mem[957] = 16'h0000;
initial mem[958] = 16'h0000;
initial mem[959] = 16'h0000;
initial mem[960] = 16'h0000;
initial mem[961] = 16'h0000;
initial mem[962] = 16'h0000;
initial mem[963] = 16'h0000;
initial mem[964] = 16'h0000;
initial mem[965] = 16'h0000;
initial mem[966] = 16'h0000;
initial mem[967] = 16'h0000;
initial mem[968] = 16'h0000;
initial mem[969] = 16'h0000;
initial mem[970] = 16'h0000;
initial mem[971] = 16'h0000;
initial mem[972] = 16'h0000;
initial mem[973] = 16'h0000;
initial mem[974] = 16'h0000;
initial mem[975] = 16'h0000;
initial mem[976] = 16'h0000;
initial mem[977] = 16'h0000;
initial mem[978] = 16'h0000;
initial mem[979] = 16'h0000;
initial mem[980] = 16'h0000;
initial mem[981] = 16'h0000;
initial mem[982] = 16'h0000;
initial mem[983] = 16'h0000;
initial mem[984] = 16'h0000;
initial mem[985] = 16'h0000;
initial mem[986] = 16'h0000;
initial mem[987] = 16'h0000;
initial mem[988] = 16'h0000;
initial mem[989] = 16'h0000;
initial mem[990] = 16'h0000;
initial mem[991] = 16'h0000;
initial mem[992] = 16'h0000;
initial mem[993] = 16'h0000;
initial mem[994] = 16'h0000;
initial mem[995] = 16'h0000;
initial mem[996] = 16'h0000;
initial mem[997] = 16'h0000;
initial mem[998] = 16'h0000;
initial mem[999] = 16'h0000;
initial mem[1000] = 16'h0000;
initial mem[1001] = 16'h0000;
initial mem[1002] = 16'h0000;
initial mem[1003] = 16'h0000;
initial mem[1004] = 16'h0000;
initial mem[1005] = 16'h0000;
initial mem[1006] = 16'h0000;
initial mem[1007] = 16'h0000;
initial mem[1008] = 16'h0000;
initial mem[1009] = 16'h0000;
initial mem[1010] = 16'h0000;
initial mem[1011] = 16'h0000;
initial mem[1012] = 16'h0000;
initial mem[1013] = 16'h0000;
initial mem[1014] = 16'h0000;
initial mem[1015] = 16'h0000;
initial mem[1016] = 16'h0000;
initial mem[1017] = 16'h0000;
initial mem[1018] = 16'h0000;
initial mem[1019] = 16'h0000;
initial mem[1020] = 16'h0000;
initial mem[1021] = 16'h0000;
initial mem[1022] = 16'h0000;
initial mem[1023] = 16'h0000;
initial mem[1024] = 16'h0000;
initial mem[1025] = 16'h0000;
initial mem[1026] = 16'h0000;
initial mem[1027] = 16'h0000;
initial mem[1028] = 16'h0000;
initial mem[1029] = 16'h0000;
initial mem[1030] = 16'h0000;
initial mem[1031] = 16'h0000;
initial mem[1032] = 16'h0000;
initial mem[1033] = 16'h0000;
initial mem[1034] = 16'h0000;
initial mem[1035] = 16'h0000;
initial mem[1036] = 16'h0000;
initial mem[1037] = 16'h0000;
initial mem[1038] = 16'h0000;
initial mem[1039] = 16'h0000;
initial mem[1040] = 16'h0000;
initial mem[1041] = 16'h0000;
initial mem[1042] = 16'h0000;
initial mem[1043] = 16'h0000;
initial mem[1044] = 16'h0000;
initial mem[1045] = 16'h0000;
initial mem[1046] = 16'h0000;
initial mem[1047] = 16'h0000;
initial mem[1048] = 16'h0000;
initial mem[1049] = 16'h0000;
initial mem[1050] = 16'h0000;
initial mem[1051] = 16'h0000;
initial mem[1052] = 16'h0000;
initial mem[1053] = 16'h0000;
initial mem[1054] = 16'h0000;
initial mem[1055] = 16'h0000;
initial mem[1056] = 16'h0000;
initial mem[1057] = 16'h0000;
initial mem[1058] = 16'h0000;
initial mem[1059] = 16'h0000;
initial mem[1060] = 16'h0000;
initial mem[1061] = 16'h0000;
initial mem[1062] = 16'h0000;
initial mem[1063] = 16'h0000;
initial mem[1064] = 16'h0000;
initial mem[1065] = 16'h0000;
initial mem[1066] = 16'h0000;
initial mem[1067] = 16'h0000;
initial mem[1068] = 16'h0000;
initial mem[1069] = 16'h0000;
initial mem[1070] = 16'h0000;
initial mem[1071] = 16'h0000;
initial mem[1072] = 16'h0000;
initial mem[1073] = 16'h0000;
initial mem[1074] = 16'h0000;
initial mem[1075] = 16'h0000;
initial mem[1076] = 16'h0000;
initial mem[1077] = 16'h0000;
initial mem[1078] = 16'h0000;
initial mem[1079] = 16'h0000;
initial mem[1080] = 16'h0000;
initial mem[1081] = 16'h0000;
initial mem[1082] = 16'h0000;
initial mem[1083] = 16'h0000;
initial mem[1084] = 16'h0000;
initial mem[1085] = 16'h0000;
initial mem[1086] = 16'h0000;
initial mem[1087] = 16'h0000;
initial mem[1088] = 16'h0000;
initial mem[1089] = 16'h0000;
initial mem[1090] = 16'h0000;
initial mem[1091] = 16'h0000;
initial mem[1092] = 16'h0000;
initial mem[1093] = 16'h0000;
initial mem[1094] = 16'h0000;
initial mem[1095] = 16'h0000;
initial mem[1096] = 16'h0000;
initial mem[1097] = 16'h0000;
initial mem[1098] = 16'h0000;
initial mem[1099] = 16'h0000;
initial mem[1100] = 16'h0000;
initial mem[1101] = 16'h0000;
initial mem[1102] = 16'h0000;
initial mem[1103] = 16'h0000;
initial mem[1104] = 16'h0000;
initial mem[1105] = 16'h0000;
initial mem[1106] = 16'h0000;
initial mem[1107] = 16'h0000;
initial mem[1108] = 16'h0000;
initial mem[1109] = 16'h0000;
initial mem[1110] = 16'h0000;
initial mem[1111] = 16'h0000;
initial mem[1112] = 16'h0000;
initial mem[1113] = 16'h0000;
initial mem[1114] = 16'h0000;
initial mem[1115] = 16'h0000;
initial mem[1116] = 16'h0000;
initial mem[1117] = 16'h0000;
initial mem[1118] = 16'h0000;
initial mem[1119] = 16'h0000;
initial mem[1120] = 16'h0000;
initial mem[1121] = 16'h0000;
initial mem[1122] = 16'h0000;
initial mem[1123] = 16'h0000;
initial mem[1124] = 16'h0000;
initial mem[1125] = 16'h0000;
initial mem[1126] = 16'h0000;
initial mem[1127] = 16'h0000;
initial mem[1128] = 16'h0000;
initial mem[1129] = 16'h0000;
initial mem[1130] = 16'h0000;
initial mem[1131] = 16'h0000;
initial mem[1132] = 16'h0000;
initial mem[1133] = 16'h0000;
initial mem[1134] = 16'h0000;
initial mem[1135] = 16'h0000;
initial mem[1136] = 16'h0000;
initial mem[1137] = 16'h0000;
initial mem[1138] = 16'h0000;
initial mem[1139] = 16'h0000;
initial mem[1140] = 16'h0000;
initial mem[1141] = 16'h0000;
initial mem[1142] = 16'h0000;
initial mem[1143] = 16'h0000;
initial mem[1144] = 16'h0000;
initial mem[1145] = 16'h0000;
initial mem[1146] = 16'h0000;
initial mem[1147] = 16'h0000;
initial mem[1148] = 16'h0000;
initial mem[1149] = 16'h0000;
initial mem[1150] = 16'h0000;
initial mem[1151] = 16'h0000;
initial mem[1152] = 16'h0000;
initial mem[1153] = 16'h0000;
initial mem[1154] = 16'h0000;
initial mem[1155] = 16'h0000;
initial mem[1156] = 16'h0000;
initial mem[1157] = 16'h0000;
initial mem[1158] = 16'h0000;
initial mem[1159] = 16'h0000;
initial mem[1160] = 16'h0000;
initial mem[1161] = 16'h0000;
initial mem[1162] = 16'h0000;
initial mem[1163] = 16'h0000;
initial mem[1164] = 16'h0000;
initial mem[1165] = 16'h0000;
initial mem[1166] = 16'h0000;
initial mem[1167] = 16'h0000;
initial mem[1168] = 16'h0000;
initial mem[1169] = 16'h0000;
initial mem[1170] = 16'h0000;
initial mem[1171] = 16'h0000;
initial mem[1172] = 16'h0000;
initial mem[1173] = 16'h0000;
initial mem[1174] = 16'h0000;
initial mem[1175] = 16'h0000;
initial mem[1176] = 16'h0000;
initial mem[1177] = 16'h0000;
initial mem[1178] = 16'h0000;
initial mem[1179] = 16'h0000;
initial mem[1180] = 16'h0000;
initial mem[1181] = 16'h0000;
initial mem[1182] = 16'h0000;
initial mem[1183] = 16'h0000;
initial mem[1184] = 16'h0000;
initial mem[1185] = 16'h0000;
initial mem[1186] = 16'h0000;
initial mem[1187] = 16'h0000;
initial mem[1188] = 16'h0000;
initial mem[1189] = 16'h0000;
initial mem[1190] = 16'h0000;
initial mem[1191] = 16'h0000;
initial mem[1192] = 16'h0000;
initial mem[1193] = 16'h0000;
initial mem[1194] = 16'h0000;
initial mem[1195] = 16'h0000;
initial mem[1196] = 16'h0000;
initial mem[1197] = 16'h0000;
initial mem[1198] = 16'h0000;
initial mem[1199] = 16'h0000;
initial mem[1200] = 16'h0000;
initial mem[1201] = 16'h0000;
initial mem[1202] = 16'h0000;
initial mem[1203] = 16'h0000;
initial mem[1204] = 16'h0000;
initial mem[1205] = 16'h0000;
initial mem[1206] = 16'h0000;
initial mem[1207] = 16'h0000;
initial mem[1208] = 16'h0000;
initial mem[1209] = 16'h0000;
initial mem[1210] = 16'h0000;
initial mem[1211] = 16'h0000;
initial mem[1212] = 16'h0000;
initial mem[1213] = 16'h0000;
initial mem[1214] = 16'h0000;
initial mem[1215] = 16'h0000;
initial mem[1216] = 16'h0000;
initial mem[1217] = 16'h0000;
initial mem[1218] = 16'h0000;
initial mem[1219] = 16'h0000;
initial mem[1220] = 16'h0000;
initial mem[1221] = 16'h0000;
initial mem[1222] = 16'h0000;
initial mem[1223] = 16'h0000;
initial mem[1224] = 16'h0000;
initial mem[1225] = 16'h0000;
initial mem[1226] = 16'h0000;
initial mem[1227] = 16'h0000;
initial mem[1228] = 16'h0000;
initial mem[1229] = 16'h0000;
initial mem[1230] = 16'h0000;
initial mem[1231] = 16'h0000;
initial mem[1232] = 16'h0000;
initial mem[1233] = 16'h0000;
initial mem[1234] = 16'h0000;
initial mem[1235] = 16'h0000;
initial mem[1236] = 16'h0000;
initial mem[1237] = 16'h0000;
initial mem[1238] = 16'h0000;
initial mem[1239] = 16'h0000;
initial mem[1240] = 16'h0000;
initial mem[1241] = 16'h0000;
initial mem[1242] = 16'h0000;
initial mem[1243] = 16'h0000;
initial mem[1244] = 16'h0000;
initial mem[1245] = 16'h0000;
initial mem[1246] = 16'h0000;
initial mem[1247] = 16'h0000;
initial mem[1248] = 16'h0000;
initial mem[1249] = 16'h0000;
initial mem[1250] = 16'h0000;
initial mem[1251] = 16'h0000;
initial mem[1252] = 16'h0000;
initial mem[1253] = 16'h0000;
initial mem[1254] = 16'h0000;
initial mem[1255] = 16'h0000;
initial mem[1256] = 16'h0000;
initial mem[1257] = 16'h0000;
initial mem[1258] = 16'h0000;
initial mem[1259] = 16'h0000;
initial mem[1260] = 16'h0000;
initial mem[1261] = 16'h0000;
initial mem[1262] = 16'h0000;
initial mem[1263] = 16'h0000;
initial mem[1264] = 16'h0000;
initial mem[1265] = 16'h0000;
initial mem[1266] = 16'h0000;
initial mem[1267] = 16'h0000;
initial mem[1268] = 16'h0000;
initial mem[1269] = 16'h0000;
initial mem[1270] = 16'h0000;
initial mem[1271] = 16'h0000;
initial mem[1272] = 16'h0000;
initial mem[1273] = 16'h0000;
initial mem[1274] = 16'h0000;
initial mem[1275] = 16'h0000;
initial mem[1276] = 16'h0000;
initial mem[1277] = 16'h0000;
initial mem[1278] = 16'h0000;
initial mem[1279] = 16'h0000;
initial mem[1280] = 16'h0000;
initial mem[1281] = 16'h0000;
initial mem[1282] = 16'h0000;
initial mem[1283] = 16'h0000;
initial mem[1284] = 16'h0000;
initial mem[1285] = 16'h0000;
initial mem[1286] = 16'h0000;
initial mem[1287] = 16'h0000;
initial mem[1288] = 16'h0000;
initial mem[1289] = 16'h0000;
initial mem[1290] = 16'h0000;
initial mem[1291] = 16'h0000;
initial mem[1292] = 16'h0000;
initial mem[1293] = 16'h0000;
initial mem[1294] = 16'h0000;
initial mem[1295] = 16'h0000;
initial mem[1296] = 16'h0000;
initial mem[1297] = 16'h0000;
initial mem[1298] = 16'h0000;
initial mem[1299] = 16'h0000;
initial mem[1300] = 16'h0000;
initial mem[1301] = 16'h0000;
initial mem[1302] = 16'h0000;
initial mem[1303] = 16'h0000;
initial mem[1304] = 16'h0000;
initial mem[1305] = 16'h0000;
initial mem[1306] = 16'h0000;
initial mem[1307] = 16'h0000;
initial mem[1308] = 16'h0000;
initial mem[1309] = 16'h0000;
initial mem[1310] = 16'h0000;
initial mem[1311] = 16'h0000;
initial mem[1312] = 16'h0000;
initial mem[1313] = 16'h0000;
initial mem[1314] = 16'h0000;
initial mem[1315] = 16'h0000;
initial mem[1316] = 16'h0000;
initial mem[1317] = 16'h0000;
initial mem[1318] = 16'h0000;
initial mem[1319] = 16'h0000;
initial mem[1320] = 16'h0000;
initial mem[1321] = 16'h0000;
initial mem[1322] = 16'h0000;
initial mem[1323] = 16'h0000;
initial mem[1324] = 16'h0000;
initial mem[1325] = 16'h0000;
initial mem[1326] = 16'h0000;
initial mem[1327] = 16'h0000;
initial mem[1328] = 16'h0000;
initial mem[1329] = 16'h0000;
initial mem[1330] = 16'h0000;
initial mem[1331] = 16'h0000;
initial mem[1332] = 16'h0000;
initial mem[1333] = 16'h0000;
initial mem[1334] = 16'h0000;
initial mem[1335] = 16'h0000;
initial mem[1336] = 16'h0000;
initial mem[1337] = 16'h0000;
initial mem[1338] = 16'h0000;
initial mem[1339] = 16'h0000;
initial mem[1340] = 16'h0000;
initial mem[1341] = 16'h0000;
initial mem[1342] = 16'h0000;
initial mem[1343] = 16'h0000;
initial mem[1344] = 16'h0000;
initial mem[1345] = 16'h0000;
initial mem[1346] = 16'h0000;
initial mem[1347] = 16'h0000;
initial mem[1348] = 16'h0000;
initial mem[1349] = 16'h0000;
initial mem[1350] = 16'h0000;
initial mem[1351] = 16'h0000;
initial mem[1352] = 16'h0000;
initial mem[1353] = 16'h0000;
initial mem[1354] = 16'h0000;
initial mem[1355] = 16'h0000;
initial mem[1356] = 16'h0000;
initial mem[1357] = 16'h0000;
initial mem[1358] = 16'h0000;
initial mem[1359] = 16'h0000;
initial mem[1360] = 16'h0000;
initial mem[1361] = 16'h0000;
initial mem[1362] = 16'h0000;
initial mem[1363] = 16'h0000;
initial mem[1364] = 16'h0000;
initial mem[1365] = 16'h0000;
initial mem[1366] = 16'h0000;
initial mem[1367] = 16'h0000;
initial mem[1368] = 16'h0000;
initial mem[1369] = 16'h0000;
initial mem[1370] = 16'h0000;
initial mem[1371] = 16'h0000;
initial mem[1372] = 16'h0000;
initial mem[1373] = 16'h0000;
initial mem[1374] = 16'h0000;
initial mem[1375] = 16'h0000;
initial mem[1376] = 16'h0000;
initial mem[1377] = 16'h0000;
initial mem[1378] = 16'h0000;
initial mem[1379] = 16'h0000;
initial mem[1380] = 16'h0000;
initial mem[1381] = 16'h0000;
initial mem[1382] = 16'h0000;
initial mem[1383] = 16'h0000;
initial mem[1384] = 16'h0000;
initial mem[1385] = 16'h0000;
initial mem[1386] = 16'h0000;
initial mem[1387] = 16'h0000;
initial mem[1388] = 16'h0000;
initial mem[1389] = 16'h0000;
initial mem[1390] = 16'h0000;
initial mem[1391] = 16'h0000;
initial mem[1392] = 16'h0000;
initial mem[1393] = 16'h0000;
initial mem[1394] = 16'h0000;
initial mem[1395] = 16'h0000;
initial mem[1396] = 16'h0000;
initial mem[1397] = 16'h0000;
initial mem[1398] = 16'h0000;
initial mem[1399] = 16'h0000;
initial mem[1400] = 16'h0000;
initial mem[1401] = 16'h0000;
initial mem[1402] = 16'h0000;
initial mem[1403] = 16'h0000;
initial mem[1404] = 16'h0000;
initial mem[1405] = 16'h0000;
initial mem[1406] = 16'h0000;
initial mem[1407] = 16'h0000;
initial mem[1408] = 16'h0000;
initial mem[1409] = 16'h0000;
initial mem[1410] = 16'h0000;
initial mem[1411] = 16'h0000;
initial mem[1412] = 16'h0000;
initial mem[1413] = 16'h0000;
initial mem[1414] = 16'h0000;
initial mem[1415] = 16'h0000;
initial mem[1416] = 16'h0000;
initial mem[1417] = 16'h0000;
initial mem[1418] = 16'h0000;
initial mem[1419] = 16'h0000;
initial mem[1420] = 16'h0000;
initial mem[1421] = 16'h0000;
initial mem[1422] = 16'h0000;
initial mem[1423] = 16'h0000;
initial mem[1424] = 16'h0000;
initial mem[1425] = 16'h0000;
initial mem[1426] = 16'h0000;
initial mem[1427] = 16'h0000;
initial mem[1428] = 16'h0000;
initial mem[1429] = 16'h0000;
initial mem[1430] = 16'h0000;
initial mem[1431] = 16'h0000;
initial mem[1432] = 16'h0000;
initial mem[1433] = 16'h0000;
initial mem[1434] = 16'h0000;
initial mem[1435] = 16'h0000;
initial mem[1436] = 16'h0000;
initial mem[1437] = 16'h0000;
initial mem[1438] = 16'h0000;
initial mem[1439] = 16'h0000;
initial mem[1440] = 16'h0000;
initial mem[1441] = 16'h0000;
initial mem[1442] = 16'h0000;
initial mem[1443] = 16'h0000;
initial mem[1444] = 16'h0000;
initial mem[1445] = 16'h0000;
initial mem[1446] = 16'h0000;
initial mem[1447] = 16'h0000;
initial mem[1448] = 16'h0000;
initial mem[1449] = 16'h0000;
initial mem[1450] = 16'h0000;
initial mem[1451] = 16'h0000;
initial mem[1452] = 16'h0000;
initial mem[1453] = 16'h0000;
initial mem[1454] = 16'h0000;
initial mem[1455] = 16'h0000;
initial mem[1456] = 16'h0000;
initial mem[1457] = 16'h0000;
initial mem[1458] = 16'h0000;
initial mem[1459] = 16'h0000;
initial mem[1460] = 16'h0000;
initial mem[1461] = 16'h0000;
initial mem[1462] = 16'h0000;
initial mem[1463] = 16'h0000;
initial mem[1464] = 16'h0000;
initial mem[1465] = 16'h0000;
initial mem[1466] = 16'h0000;
initial mem[1467] = 16'h0000;
initial mem[1468] = 16'h0000;
initial mem[1469] = 16'h0000;
initial mem[1470] = 16'h0000;
initial mem[1471] = 16'h0000;
initial mem[1472] = 16'h0000;
initial mem[1473] = 16'h0000;
initial mem[1474] = 16'h0000;
initial mem[1475] = 16'h0000;
initial mem[1476] = 16'h0000;
initial mem[1477] = 16'h0000;
initial mem[1478] = 16'h0000;
initial mem[1479] = 16'h0000;
initial mem[1480] = 16'h0000;
initial mem[1481] = 16'h0000;
initial mem[1482] = 16'h0000;
initial mem[1483] = 16'h0000;
initial mem[1484] = 16'h0000;
initial mem[1485] = 16'h0000;
initial mem[1486] = 16'h0000;
initial mem[1487] = 16'h0000;
initial mem[1488] = 16'h0000;
initial mem[1489] = 16'h0000;
initial mem[1490] = 16'h0000;
initial mem[1491] = 16'h0000;
initial mem[1492] = 16'h0000;
initial mem[1493] = 16'h0000;
initial mem[1494] = 16'h0000;
initial mem[1495] = 16'h0000;
initial mem[1496] = 16'h0000;
initial mem[1497] = 16'h0000;
initial mem[1498] = 16'h0000;
initial mem[1499] = 16'h0000;
initial mem[1500] = 16'h0000;
initial mem[1501] = 16'h0000;
initial mem[1502] = 16'h0000;
initial mem[1503] = 16'h0000;
initial mem[1504] = 16'h0000;
initial mem[1505] = 16'h0000;
initial mem[1506] = 16'h0000;
initial mem[1507] = 16'h0000;
initial mem[1508] = 16'h0000;
initial mem[1509] = 16'h0000;
initial mem[1510] = 16'h0000;
initial mem[1511] = 16'h0000;
initial mem[1512] = 16'h0000;
initial mem[1513] = 16'h0000;
initial mem[1514] = 16'h0000;
initial mem[1515] = 16'h0000;
initial mem[1516] = 16'h0000;
initial mem[1517] = 16'h0000;
initial mem[1518] = 16'h0000;
initial mem[1519] = 16'h0000;
initial mem[1520] = 16'h0000;
initial mem[1521] = 16'h0000;
initial mem[1522] = 16'h0000;
initial mem[1523] = 16'h0000;
initial mem[1524] = 16'h0000;
initial mem[1525] = 16'h0000;
initial mem[1526] = 16'h0000;
initial mem[1527] = 16'h0000;
initial mem[1528] = 16'h0000;
initial mem[1529] = 16'h0000;
initial mem[1530] = 16'h0000;
initial mem[1531] = 16'h0000;
initial mem[1532] = 16'h0000;
initial mem[1533] = 16'h0000;
initial mem[1534] = 16'h0000;
initial mem[1535] = 16'h0000;
initial mem[1536] = 16'h0000;
initial mem[1537] = 16'h0000;
initial mem[1538] = 16'h0000;
initial mem[1539] = 16'h0000;
initial mem[1540] = 16'h0000;
initial mem[1541] = 16'h0000;
initial mem[1542] = 16'h0000;
initial mem[1543] = 16'h0000;
initial mem[1544] = 16'h0000;
initial mem[1545] = 16'h0000;
initial mem[1546] = 16'h0000;
initial mem[1547] = 16'h0000;
initial mem[1548] = 16'h0000;
initial mem[1549] = 16'h0000;
initial mem[1550] = 16'h0000;
initial mem[1551] = 16'h0000;
initial mem[1552] = 16'h0000;
initial mem[1553] = 16'h0000;
initial mem[1554] = 16'h0000;
initial mem[1555] = 16'h0000;
initial mem[1556] = 16'h0000;
initial mem[1557] = 16'h0000;
initial mem[1558] = 16'h0000;
initial mem[1559] = 16'h0000;
initial mem[1560] = 16'h0000;
initial mem[1561] = 16'h0000;
initial mem[1562] = 16'h0000;
initial mem[1563] = 16'h0000;
initial mem[1564] = 16'h0000;
initial mem[1565] = 16'h0000;
initial mem[1566] = 16'h0000;
initial mem[1567] = 16'h0000;
initial mem[1568] = 16'h0000;
initial mem[1569] = 16'h0000;
initial mem[1570] = 16'h0000;
initial mem[1571] = 16'h0000;
initial mem[1572] = 16'h0000;
initial mem[1573] = 16'h0000;
initial mem[1574] = 16'h0000;
initial mem[1575] = 16'h0000;
initial mem[1576] = 16'h0000;
initial mem[1577] = 16'h0000;
initial mem[1578] = 16'h0000;
initial mem[1579] = 16'h0000;
initial mem[1580] = 16'h0000;
initial mem[1581] = 16'h0000;
initial mem[1582] = 16'h0000;
initial mem[1583] = 16'h0000;
initial mem[1584] = 16'h0000;
initial mem[1585] = 16'h0000;
initial mem[1586] = 16'h0000;
initial mem[1587] = 16'h0000;
initial mem[1588] = 16'h0000;
initial mem[1589] = 16'h0000;
initial mem[1590] = 16'h0000;
initial mem[1591] = 16'h0000;
initial mem[1592] = 16'h0000;
initial mem[1593] = 16'h0000;
initial mem[1594] = 16'h0000;
initial mem[1595] = 16'h0000;
initial mem[1596] = 16'h0000;
initial mem[1597] = 16'h0000;
initial mem[1598] = 16'h0000;
initial mem[1599] = 16'h0000;
initial mem[1600] = 16'h0000;
initial mem[1601] = 16'h0000;
initial mem[1602] = 16'h0000;
initial mem[1603] = 16'h0000;
initial mem[1604] = 16'h0000;
initial mem[1605] = 16'h0000;
initial mem[1606] = 16'h0000;
initial mem[1607] = 16'h0000;
initial mem[1608] = 16'h0000;
initial mem[1609] = 16'h0000;
initial mem[1610] = 16'h0000;
initial mem[1611] = 16'h0000;
initial mem[1612] = 16'h0000;
initial mem[1613] = 16'h0000;
initial mem[1614] = 16'h0000;
initial mem[1615] = 16'h0000;
initial mem[1616] = 16'h0000;
initial mem[1617] = 16'h0000;
initial mem[1618] = 16'h0000;
initial mem[1619] = 16'h0000;
initial mem[1620] = 16'h0000;
initial mem[1621] = 16'h0000;
initial mem[1622] = 16'h0000;
initial mem[1623] = 16'h0000;
initial mem[1624] = 16'h0000;
initial mem[1625] = 16'h0000;
initial mem[1626] = 16'h0000;
initial mem[1627] = 16'h0000;
initial mem[1628] = 16'h0000;
initial mem[1629] = 16'h0000;
initial mem[1630] = 16'h0000;
initial mem[1631] = 16'h0000;
initial mem[1632] = 16'h0000;
initial mem[1633] = 16'h0000;
initial mem[1634] = 16'h0000;
initial mem[1635] = 16'h0000;
initial mem[1636] = 16'h0000;
initial mem[1637] = 16'h0000;
initial mem[1638] = 16'h0000;
initial mem[1639] = 16'h0000;
initial mem[1640] = 16'h0000;
initial mem[1641] = 16'h0000;
initial mem[1642] = 16'h0000;
initial mem[1643] = 16'h0000;
initial mem[1644] = 16'h0000;
initial mem[1645] = 16'h0000;
initial mem[1646] = 16'h0000;
initial mem[1647] = 16'h0000;
initial mem[1648] = 16'h0000;
initial mem[1649] = 16'h0000;
initial mem[1650] = 16'h0000;
initial mem[1651] = 16'h0000;
initial mem[1652] = 16'h0000;
initial mem[1653] = 16'h0000;
initial mem[1654] = 16'h0000;
initial mem[1655] = 16'h0000;
initial mem[1656] = 16'h0000;
initial mem[1657] = 16'h0000;
initial mem[1658] = 16'h0000;
initial mem[1659] = 16'h0000;
initial mem[1660] = 16'h0000;
initial mem[1661] = 16'h0000;
initial mem[1662] = 16'h0000;
initial mem[1663] = 16'h0000;
initial mem[1664] = 16'h0000;
initial mem[1665] = 16'h0000;
initial mem[1666] = 16'h0000;
initial mem[1667] = 16'h0000;
initial mem[1668] = 16'h0000;
initial mem[1669] = 16'h0000;
initial mem[1670] = 16'h0000;
initial mem[1671] = 16'h0000;
initial mem[1672] = 16'h0000;
initial mem[1673] = 16'h0000;
initial mem[1674] = 16'h0000;
initial mem[1675] = 16'h0000;
initial mem[1676] = 16'h0000;
initial mem[1677] = 16'h0000;
initial mem[1678] = 16'h0000;
initial mem[1679] = 16'h0000;
initial mem[1680] = 16'h0000;
initial mem[1681] = 16'h0000;
initial mem[1682] = 16'h0000;
initial mem[1683] = 16'h0000;
initial mem[1684] = 16'h0000;
initial mem[1685] = 16'h0000;
initial mem[1686] = 16'h0000;
initial mem[1687] = 16'h0000;
initial mem[1688] = 16'h0000;
initial mem[1689] = 16'h0000;
initial mem[1690] = 16'h0000;
initial mem[1691] = 16'h0000;
initial mem[1692] = 16'h0000;
initial mem[1693] = 16'h0000;
initial mem[1694] = 16'h0000;
initial mem[1695] = 16'h0000;
initial mem[1696] = 16'h0000;
initial mem[1697] = 16'h0000;
initial mem[1698] = 16'h0000;
initial mem[1699] = 16'h0000;
initial mem[1700] = 16'h0000;
initial mem[1701] = 16'h0000;
initial mem[1702] = 16'h0000;
initial mem[1703] = 16'h0000;
initial mem[1704] = 16'h0000;
initial mem[1705] = 16'h0000;
initial mem[1706] = 16'h0000;
initial mem[1707] = 16'h0000;
initial mem[1708] = 16'h0000;
initial mem[1709] = 16'h0000;
initial mem[1710] = 16'h0000;
initial mem[1711] = 16'h0000;
initial mem[1712] = 16'h0000;
initial mem[1713] = 16'h0000;
initial mem[1714] = 16'h0000;
initial mem[1715] = 16'h0000;
initial mem[1716] = 16'h0000;
initial mem[1717] = 16'h0000;
initial mem[1718] = 16'h0000;
initial mem[1719] = 16'h0000;
initial mem[1720] = 16'h0000;
initial mem[1721] = 16'h0000;
initial mem[1722] = 16'h0000;
initial mem[1723] = 16'h0000;
initial mem[1724] = 16'h0000;
initial mem[1725] = 16'h0000;
initial mem[1726] = 16'h0000;
initial mem[1727] = 16'h0000;
initial mem[1728] = 16'h0000;
initial mem[1729] = 16'h0000;
initial mem[1730] = 16'h0000;
initial mem[1731] = 16'h0000;
initial mem[1732] = 16'h0000;
initial mem[1733] = 16'h0000;
initial mem[1734] = 16'h0000;
initial mem[1735] = 16'h0000;
initial mem[1736] = 16'h0000;
initial mem[1737] = 16'h0000;
initial mem[1738] = 16'h0000;
initial mem[1739] = 16'h0000;
initial mem[1740] = 16'h0000;
initial mem[1741] = 16'h0000;
initial mem[1742] = 16'h0000;
initial mem[1743] = 16'h0000;
initial mem[1744] = 16'h0000;
initial mem[1745] = 16'h0000;
initial mem[1746] = 16'h0000;
initial mem[1747] = 16'h0000;
initial mem[1748] = 16'h0000;
initial mem[1749] = 16'h0000;
initial mem[1750] = 16'h0000;
initial mem[1751] = 16'h0000;
initial mem[1752] = 16'h0000;
initial mem[1753] = 16'h0000;
initial mem[1754] = 16'h0000;
initial mem[1755] = 16'h0000;
initial mem[1756] = 16'h0000;
initial mem[1757] = 16'h0000;
initial mem[1758] = 16'h0000;
initial mem[1759] = 16'h0000;
initial mem[1760] = 16'h0000;
initial mem[1761] = 16'h0000;
initial mem[1762] = 16'h0000;
initial mem[1763] = 16'h0000;
initial mem[1764] = 16'h0000;
initial mem[1765] = 16'h0000;
initial mem[1766] = 16'h0000;
initial mem[1767] = 16'h0000;
initial mem[1768] = 16'h0000;
initial mem[1769] = 16'h0000;
initial mem[1770] = 16'h0000;
initial mem[1771] = 16'h0000;
initial mem[1772] = 16'h0000;
initial mem[1773] = 16'h0000;
initial mem[1774] = 16'h0000;
initial mem[1775] = 16'h0000;
initial mem[1776] = 16'h0000;
initial mem[1777] = 16'h0000;
initial mem[1778] = 16'h0000;
initial mem[1779] = 16'h0000;
initial mem[1780] = 16'h0000;
initial mem[1781] = 16'h0000;
initial mem[1782] = 16'h0000;
initial mem[1783] = 16'h0000;
initial mem[1784] = 16'h0000;
initial mem[1785] = 16'h0000;
initial mem[1786] = 16'h0000;
initial mem[1787] = 16'h0000;
initial mem[1788] = 16'h0000;
initial mem[1789] = 16'h0000;
initial mem[1790] = 16'h0000;
initial mem[1791] = 16'h0000;
initial mem[1792] = 16'h0000;
initial mem[1793] = 16'h0000;
initial mem[1794] = 16'h0000;
initial mem[1795] = 16'h0000;
initial mem[1796] = 16'h0000;
initial mem[1797] = 16'h0000;
initial mem[1798] = 16'h0000;
initial mem[1799] = 16'h0000;
initial mem[1800] = 16'h0000;
initial mem[1801] = 16'h0000;
initial mem[1802] = 16'h0000;
initial mem[1803] = 16'h0000;
initial mem[1804] = 16'h0000;
initial mem[1805] = 16'h0000;
initial mem[1806] = 16'h0000;
initial mem[1807] = 16'h0000;
initial mem[1808] = 16'h0000;
initial mem[1809] = 16'h0000;
initial mem[1810] = 16'h0000;
initial mem[1811] = 16'h0000;
initial mem[1812] = 16'h0000;
initial mem[1813] = 16'h0000;
initial mem[1814] = 16'h0000;
initial mem[1815] = 16'h0000;
initial mem[1816] = 16'h0000;
initial mem[1817] = 16'h0000;
initial mem[1818] = 16'h0000;
initial mem[1819] = 16'h0000;
initial mem[1820] = 16'h0000;
initial mem[1821] = 16'h0000;
initial mem[1822] = 16'h0000;
initial mem[1823] = 16'h0000;
initial mem[1824] = 16'h0000;
initial mem[1825] = 16'h0000;
initial mem[1826] = 16'h0000;
initial mem[1827] = 16'h0000;
initial mem[1828] = 16'h0000;
initial mem[1829] = 16'h0000;
initial mem[1830] = 16'h0000;
initial mem[1831] = 16'h0000;
initial mem[1832] = 16'h0000;
initial mem[1833] = 16'h0000;
initial mem[1834] = 16'h0000;
initial mem[1835] = 16'h0000;
initial mem[1836] = 16'h0000;
initial mem[1837] = 16'h0000;
initial mem[1838] = 16'h0000;
initial mem[1839] = 16'h0000;
initial mem[1840] = 16'h0000;
initial mem[1841] = 16'h0000;
initial mem[1842] = 16'h0000;
initial mem[1843] = 16'h0000;
initial mem[1844] = 16'h0000;
initial mem[1845] = 16'h0000;
initial mem[1846] = 16'h0000;
initial mem[1847] = 16'h0000;
initial mem[1848] = 16'h0000;
initial mem[1849] = 16'h0000;
initial mem[1850] = 16'h0000;
initial mem[1851] = 16'h0000;
initial mem[1852] = 16'h0000;
initial mem[1853] = 16'h0000;
initial mem[1854] = 16'h0000;
initial mem[1855] = 16'h0000;
initial mem[1856] = 16'h0000;
initial mem[1857] = 16'h0000;
initial mem[1858] = 16'h0000;
initial mem[1859] = 16'h0000;
initial mem[1860] = 16'h0000;
initial mem[1861] = 16'h0000;
initial mem[1862] = 16'h0000;
initial mem[1863] = 16'h0000;
initial mem[1864] = 16'h0000;
initial mem[1865] = 16'h0000;
initial mem[1866] = 16'h0000;
initial mem[1867] = 16'h0000;
initial mem[1868] = 16'h0000;
initial mem[1869] = 16'h0000;
initial mem[1870] = 16'h0000;
initial mem[1871] = 16'h0000;
initial mem[1872] = 16'h0000;
initial mem[1873] = 16'h0000;
initial mem[1874] = 16'h0000;
initial mem[1875] = 16'h0000;
initial mem[1876] = 16'h0000;
initial mem[1877] = 16'h0000;
initial mem[1878] = 16'h0000;
initial mem[1879] = 16'h0000;
initial mem[1880] = 16'h0000;
initial mem[1881] = 16'h0000;
initial mem[1882] = 16'h0000;
initial mem[1883] = 16'h0000;
initial mem[1884] = 16'h0000;
initial mem[1885] = 16'h0000;
initial mem[1886] = 16'h0000;
initial mem[1887] = 16'h0000;
initial mem[1888] = 16'h0000;
initial mem[1889] = 16'h0000;
initial mem[1890] = 16'h0000;
initial mem[1891] = 16'h0000;
initial mem[1892] = 16'h0000;
initial mem[1893] = 16'h0000;
initial mem[1894] = 16'h0000;
initial mem[1895] = 16'h0000;
initial mem[1896] = 16'h0000;
initial mem[1897] = 16'h0000;
initial mem[1898] = 16'h0000;
initial mem[1899] = 16'h0000;
initial mem[1900] = 16'h0000;
initial mem[1901] = 16'h0000;
initial mem[1902] = 16'h0000;
initial mem[1903] = 16'h0000;
initial mem[1904] = 16'h0000;
initial mem[1905] = 16'h0000;
initial mem[1906] = 16'h0000;
initial mem[1907] = 16'h0000;
initial mem[1908] = 16'h0000;
initial mem[1909] = 16'h0000;
initial mem[1910] = 16'h0000;
initial mem[1911] = 16'h0000;
initial mem[1912] = 16'h0000;
initial mem[1913] = 16'h0000;
initial mem[1914] = 16'h0000;
initial mem[1915] = 16'h0000;
initial mem[1916] = 16'h0000;
initial mem[1917] = 16'h0000;
initial mem[1918] = 16'h0000;
initial mem[1919] = 16'h0000;
initial mem[1920] = 16'h0000;
initial mem[1921] = 16'h0000;
initial mem[1922] = 16'h0000;
initial mem[1923] = 16'h0000;
initial mem[1924] = 16'h0000;
initial mem[1925] = 16'h0000;
initial mem[1926] = 16'h0000;
initial mem[1927] = 16'h0000;
initial mem[1928] = 16'h0000;
initial mem[1929] = 16'h0000;
initial mem[1930] = 16'h0000;
initial mem[1931] = 16'h0000;
initial mem[1932] = 16'h0000;
initial mem[1933] = 16'h0000;
initial mem[1934] = 16'h0000;
initial mem[1935] = 16'h0000;
initial mem[1936] = 16'h0000;
initial mem[1937] = 16'h0000;
initial mem[1938] = 16'h0000;
initial mem[1939] = 16'h0000;
initial mem[1940] = 16'h0000;
initial mem[1941] = 16'h0000;
initial mem[1942] = 16'h0000;
initial mem[1943] = 16'h0000;
initial mem[1944] = 16'h0000;
initial mem[1945] = 16'h0000;
initial mem[1946] = 16'h0000;
initial mem[1947] = 16'h0000;
initial mem[1948] = 16'h0000;
initial mem[1949] = 16'h0000;
initial mem[1950] = 16'h0000;
initial mem[1951] = 16'h0000;
initial mem[1952] = 16'h0000;
initial mem[1953] = 16'h0000;
initial mem[1954] = 16'h0000;
initial mem[1955] = 16'h0000;
initial mem[1956] = 16'h0000;
initial mem[1957] = 16'h0000;
initial mem[1958] = 16'h0000;
initial mem[1959] = 16'h0000;
initial mem[1960] = 16'h0000;
initial mem[1961] = 16'h0000;
initial mem[1962] = 16'h0000;
initial mem[1963] = 16'h0000;
initial mem[1964] = 16'h0000;
initial mem[1965] = 16'h0000;
initial mem[1966] = 16'h0000;
initial mem[1967] = 16'h0000;
initial mem[1968] = 16'h0000;
initial mem[1969] = 16'h0000;
initial mem[1970] = 16'h0000;
initial mem[1971] = 16'h0000;
initial mem[1972] = 16'h0000;
initial mem[1973] = 16'h0000;
initial mem[1974] = 16'h0000;
initial mem[1975] = 16'h0000;
initial mem[1976] = 16'h0000;
initial mem[1977] = 16'h0000;
initial mem[1978] = 16'h0000;
initial mem[1979] = 16'h0000;
initial mem[1980] = 16'h0000;
initial mem[1981] = 16'h0000;
initial mem[1982] = 16'h0000;
initial mem[1983] = 16'h0000;
initial mem[1984] = 16'h0000;
initial mem[1985] = 16'h0000;
initial mem[1986] = 16'h0000;
initial mem[1987] = 16'h0000;
initial mem[1988] = 16'h0000;
initial mem[1989] = 16'h0000;
initial mem[1990] = 16'h0000;
initial mem[1991] = 16'h0000;
initial mem[1992] = 16'h0000;
initial mem[1993] = 16'h0000;
initial mem[1994] = 16'h0000;
initial mem[1995] = 16'h0000;
initial mem[1996] = 16'h0000;
initial mem[1997] = 16'h0000;
initial mem[1998] = 16'h0000;
initial mem[1999] = 16'h0000;
initial mem[2000] = 16'h0000;
initial mem[2001] = 16'h0000;
initial mem[2002] = 16'h0000;
initial mem[2003] = 16'h0000;
initial mem[2004] = 16'h0000;
initial mem[2005] = 16'h0000;
initial mem[2006] = 16'h0000;
initial mem[2007] = 16'h0000;
initial mem[2008] = 16'h0000;
initial mem[2009] = 16'h0000;
initial mem[2010] = 16'h0000;
initial mem[2011] = 16'h0000;
initial mem[2012] = 16'h0000;
initial mem[2013] = 16'h0000;
initial mem[2014] = 16'h0000;
initial mem[2015] = 16'h0000;
initial mem[2016] = 16'h0000;
initial mem[2017] = 16'h0000;
initial mem[2018] = 16'h0000;
initial mem[2019] = 16'h0000;
initial mem[2020] = 16'h0000;
initial mem[2021] = 16'h0000;
initial mem[2022] = 16'h0000;
initial mem[2023] = 16'h0000;
initial mem[2024] = 16'h0000;
initial mem[2025] = 16'h0000;
initial mem[2026] = 16'h0000;
initial mem[2027] = 16'h0000;
initial mem[2028] = 16'h0000;
initial mem[2029] = 16'h0000;
initial mem[2030] = 16'h0000;
initial mem[2031] = 16'h0000;
initial mem[2032] = 16'h0000;
initial mem[2033] = 16'h0000;
initial mem[2034] = 16'h0000;
initial mem[2035] = 16'h0000;
initial mem[2036] = 16'h0000;
initial mem[2037] = 16'h0000;
initial mem[2038] = 16'h0000;
initial mem[2039] = 16'h0000;
initial mem[2040] = 16'h0000;
initial mem[2041] = 16'h0000;
initial mem[2042] = 16'h0000;
initial mem[2043] = 16'h0000;
initial mem[2044] = 16'h0000;
initial mem[2045] = 16'h0000;
initial mem[2046] = 16'h0000;
initial mem[2047] = 16'h0000;
initial mem[2048] = 16'h0000;
initial mem[2049] = 16'h0000;
initial mem[2050] = 16'h0000;
initial mem[2051] = 16'h0000;
initial mem[2052] = 16'h0000;
initial mem[2053] = 16'h0000;
initial mem[2054] = 16'h0000;
initial mem[2055] = 16'h0000;
initial mem[2056] = 16'h0000;
initial mem[2057] = 16'h0000;
initial mem[2058] = 16'h0000;
initial mem[2059] = 16'h0000;
initial mem[2060] = 16'h0000;
initial mem[2061] = 16'h0000;
initial mem[2062] = 16'h0000;
initial mem[2063] = 16'h0000;
initial mem[2064] = 16'h0000;
initial mem[2065] = 16'h0000;
initial mem[2066] = 16'h0000;
initial mem[2067] = 16'h0000;
initial mem[2068] = 16'h0000;
initial mem[2069] = 16'h0000;
initial mem[2070] = 16'h0000;
initial mem[2071] = 16'h0000;
initial mem[2072] = 16'h0000;
initial mem[2073] = 16'h0000;
initial mem[2074] = 16'h0000;
initial mem[2075] = 16'h0000;
initial mem[2076] = 16'h0000;
initial mem[2077] = 16'h0000;
initial mem[2078] = 16'h0000;
initial mem[2079] = 16'h0000;
initial mem[2080] = 16'h0000;
initial mem[2081] = 16'h0000;
initial mem[2082] = 16'h0000;
initial mem[2083] = 16'h0000;
initial mem[2084] = 16'h0000;
initial mem[2085] = 16'h0000;
initial mem[2086] = 16'h0000;
initial mem[2087] = 16'h0000;
initial mem[2088] = 16'h0000;
initial mem[2089] = 16'h0000;
initial mem[2090] = 16'h0000;
initial mem[2091] = 16'h0000;
initial mem[2092] = 16'h0000;
initial mem[2093] = 16'h0000;
initial mem[2094] = 16'h0000;
initial mem[2095] = 16'h0000;
initial mem[2096] = 16'h0000;
initial mem[2097] = 16'h0000;
initial mem[2098] = 16'h0000;
initial mem[2099] = 16'h0000;
initial mem[2100] = 16'h0000;
initial mem[2101] = 16'h0000;
initial mem[2102] = 16'h0000;
initial mem[2103] = 16'h0000;
initial mem[2104] = 16'h0000;
initial mem[2105] = 16'h0000;
initial mem[2106] = 16'h0000;
initial mem[2107] = 16'h0000;
initial mem[2108] = 16'h0000;
initial mem[2109] = 16'h0000;
initial mem[2110] = 16'h0000;
initial mem[2111] = 16'h0000;
initial mem[2112] = 16'h0000;
initial mem[2113] = 16'h0000;
initial mem[2114] = 16'h0000;
initial mem[2115] = 16'h0000;
initial mem[2116] = 16'h0000;
initial mem[2117] = 16'h0000;
initial mem[2118] = 16'h0000;
initial mem[2119] = 16'h0000;
initial mem[2120] = 16'h0000;
initial mem[2121] = 16'h0000;
initial mem[2122] = 16'h0000;
initial mem[2123] = 16'h0000;
initial mem[2124] = 16'h0000;
initial mem[2125] = 16'h0000;
initial mem[2126] = 16'h0000;
initial mem[2127] = 16'h0000;
initial mem[2128] = 16'h0000;
initial mem[2129] = 16'h0000;
initial mem[2130] = 16'h0000;
initial mem[2131] = 16'h0000;
initial mem[2132] = 16'h0000;
initial mem[2133] = 16'h0000;
initial mem[2134] = 16'h0000;
initial mem[2135] = 16'h0000;
initial mem[2136] = 16'h0000;
initial mem[2137] = 16'h0000;
initial mem[2138] = 16'h0000;
initial mem[2139] = 16'h0000;
initial mem[2140] = 16'h0000;
initial mem[2141] = 16'h0000;
initial mem[2142] = 16'h0000;
initial mem[2143] = 16'h0000;
initial mem[2144] = 16'h0000;
initial mem[2145] = 16'h0000;
initial mem[2146] = 16'h0000;
initial mem[2147] = 16'h0000;
initial mem[2148] = 16'h0000;
initial mem[2149] = 16'h0000;
initial mem[2150] = 16'h0000;
initial mem[2151] = 16'h0000;
initial mem[2152] = 16'h0000;
initial mem[2153] = 16'h0000;
initial mem[2154] = 16'h0000;
initial mem[2155] = 16'h0000;
initial mem[2156] = 16'h0000;
initial mem[2157] = 16'h0000;
initial mem[2158] = 16'h0000;
initial mem[2159] = 16'h0000;
initial mem[2160] = 16'h0000;
initial mem[2161] = 16'h0000;
initial mem[2162] = 16'h0000;
initial mem[2163] = 16'h0000;
initial mem[2164] = 16'h0000;
initial mem[2165] = 16'h0000;
initial mem[2166] = 16'h0000;
initial mem[2167] = 16'h0000;
initial mem[2168] = 16'h0000;
initial mem[2169] = 16'h0000;
initial mem[2170] = 16'h0000;
initial mem[2171] = 16'h0000;
initial mem[2172] = 16'h0000;
initial mem[2173] = 16'h0000;
initial mem[2174] = 16'h0000;
initial mem[2175] = 16'h0000;
initial mem[2176] = 16'h0000;
initial mem[2177] = 16'h0000;
initial mem[2178] = 16'h0000;
initial mem[2179] = 16'h0000;
initial mem[2180] = 16'h0000;
initial mem[2181] = 16'h0000;
initial mem[2182] = 16'h0000;
initial mem[2183] = 16'h0000;
initial mem[2184] = 16'h0000;
initial mem[2185] = 16'h0000;
initial mem[2186] = 16'h0000;
initial mem[2187] = 16'h0000;
initial mem[2188] = 16'h0000;
initial mem[2189] = 16'h0000;
initial mem[2190] = 16'h0000;
initial mem[2191] = 16'h0000;
initial mem[2192] = 16'h0000;
initial mem[2193] = 16'h0000;
initial mem[2194] = 16'h0000;
initial mem[2195] = 16'h0000;
initial mem[2196] = 16'h0000;
initial mem[2197] = 16'h0000;
initial mem[2198] = 16'h0000;
initial mem[2199] = 16'h0000;
initial mem[2200] = 16'h0000;
initial mem[2201] = 16'h0000;
initial mem[2202] = 16'h0000;
initial mem[2203] = 16'h0000;
initial mem[2204] = 16'h0000;
initial mem[2205] = 16'h0000;
initial mem[2206] = 16'h0000;
initial mem[2207] = 16'h0000;
initial mem[2208] = 16'h0000;
initial mem[2209] = 16'h0000;
initial mem[2210] = 16'h0000;
initial mem[2211] = 16'h0000;
initial mem[2212] = 16'h0000;
initial mem[2213] = 16'h0000;
initial mem[2214] = 16'h0000;
initial mem[2215] = 16'h0000;
initial mem[2216] = 16'h0000;
initial mem[2217] = 16'h0000;
initial mem[2218] = 16'h0000;
initial mem[2219] = 16'h0000;
initial mem[2220] = 16'h0000;
initial mem[2221] = 16'h0000;
initial mem[2222] = 16'h0000;
initial mem[2223] = 16'h0000;
initial mem[2224] = 16'h0000;
initial mem[2225] = 16'h0000;
initial mem[2226] = 16'h0000;
initial mem[2227] = 16'h0000;
initial mem[2228] = 16'h0000;
initial mem[2229] = 16'h0000;
initial mem[2230] = 16'h0000;
initial mem[2231] = 16'h0000;
initial mem[2232] = 16'h0000;
initial mem[2233] = 16'h0000;
initial mem[2234] = 16'h0000;
initial mem[2235] = 16'h0000;
initial mem[2236] = 16'h0000;
initial mem[2237] = 16'h0000;
initial mem[2238] = 16'h0000;
initial mem[2239] = 16'h0000;
initial mem[2240] = 16'h0000;
initial mem[2241] = 16'h0000;
initial mem[2242] = 16'h0000;
initial mem[2243] = 16'h0000;
initial mem[2244] = 16'h0000;
initial mem[2245] = 16'h0000;
initial mem[2246] = 16'h0000;
initial mem[2247] = 16'h0000;
initial mem[2248] = 16'h0000;
initial mem[2249] = 16'h0000;
initial mem[2250] = 16'h0000;
initial mem[2251] = 16'h0000;
initial mem[2252] = 16'h0000;
initial mem[2253] = 16'h0000;
initial mem[2254] = 16'h0000;
initial mem[2255] = 16'h0000;
initial mem[2256] = 16'h0000;
initial mem[2257] = 16'h0000;
initial mem[2258] = 16'h0000;
initial mem[2259] = 16'h0000;
initial mem[2260] = 16'h0000;
initial mem[2261] = 16'h0000;
initial mem[2262] = 16'h0000;
initial mem[2263] = 16'h0000;
initial mem[2264] = 16'h0000;
initial mem[2265] = 16'h0000;
initial mem[2266] = 16'h0000;
initial mem[2267] = 16'h0000;
initial mem[2268] = 16'h0000;
initial mem[2269] = 16'h0000;
initial mem[2270] = 16'h0000;
initial mem[2271] = 16'h0000;
initial mem[2272] = 16'h0000;
initial mem[2273] = 16'h0000;
initial mem[2274] = 16'h0000;
initial mem[2275] = 16'h0000;
initial mem[2276] = 16'h0000;
initial mem[2277] = 16'h0000;
initial mem[2278] = 16'h0000;
initial mem[2279] = 16'h0000;
initial mem[2280] = 16'h0000;
initial mem[2281] = 16'h0000;
initial mem[2282] = 16'h0000;
initial mem[2283] = 16'h0000;
initial mem[2284] = 16'h0000;
initial mem[2285] = 16'h0000;
initial mem[2286] = 16'h0000;
initial mem[2287] = 16'h0000;
initial mem[2288] = 16'h0000;
initial mem[2289] = 16'h0000;
initial mem[2290] = 16'h0000;
initial mem[2291] = 16'h0000;
initial mem[2292] = 16'h0000;
initial mem[2293] = 16'h0000;
initial mem[2294] = 16'h0000;
initial mem[2295] = 16'h0000;
initial mem[2296] = 16'h0000;
initial mem[2297] = 16'h0000;
initial mem[2298] = 16'h0000;
initial mem[2299] = 16'h0000;
initial mem[2300] = 16'h0000;
initial mem[2301] = 16'h0000;
initial mem[2302] = 16'h0000;
initial mem[2303] = 16'h0000;
initial mem[2304] = 16'h0000;
initial mem[2305] = 16'h0000;
initial mem[2306] = 16'h0000;
initial mem[2307] = 16'h0000;
initial mem[2308] = 16'h0000;
initial mem[2309] = 16'h0000;
initial mem[2310] = 16'h0000;
initial mem[2311] = 16'h0000;
initial mem[2312] = 16'h0000;
initial mem[2313] = 16'h0000;
initial mem[2314] = 16'h0000;
initial mem[2315] = 16'h0000;
initial mem[2316] = 16'h0000;
initial mem[2317] = 16'h0000;
initial mem[2318] = 16'h0000;
initial mem[2319] = 16'h0000;
initial mem[2320] = 16'h0000;
initial mem[2321] = 16'h0000;
initial mem[2322] = 16'h0000;
initial mem[2323] = 16'h0000;
initial mem[2324] = 16'h0000;
initial mem[2325] = 16'h0000;
initial mem[2326] = 16'h0000;
initial mem[2327] = 16'h0000;
initial mem[2328] = 16'h0000;
initial mem[2329] = 16'h0000;
initial mem[2330] = 16'h0000;
initial mem[2331] = 16'h0000;
initial mem[2332] = 16'h0000;
initial mem[2333] = 16'h0000;
initial mem[2334] = 16'h0000;
initial mem[2335] = 16'h0000;
initial mem[2336] = 16'h0000;
initial mem[2337] = 16'h0000;
initial mem[2338] = 16'h0000;
initial mem[2339] = 16'h0000;
initial mem[2340] = 16'h0000;
initial mem[2341] = 16'h0000;
initial mem[2342] = 16'h0000;
initial mem[2343] = 16'h0000;
initial mem[2344] = 16'h0000;
initial mem[2345] = 16'h0000;
initial mem[2346] = 16'h0000;
initial mem[2347] = 16'h0000;
initial mem[2348] = 16'h0000;
initial mem[2349] = 16'h0000;
initial mem[2350] = 16'h0000;
initial mem[2351] = 16'h0000;
initial mem[2352] = 16'h0000;
initial mem[2353] = 16'h0000;
initial mem[2354] = 16'h0000;
initial mem[2355] = 16'h0000;
initial mem[2356] = 16'h0000;
initial mem[2357] = 16'h0000;
initial mem[2358] = 16'h0000;
initial mem[2359] = 16'h0000;
initial mem[2360] = 16'h0000;
initial mem[2361] = 16'h0000;
initial mem[2362] = 16'h0000;
initial mem[2363] = 16'h0000;
initial mem[2364] = 16'h0000;
initial mem[2365] = 16'h0000;
initial mem[2366] = 16'h0000;
initial mem[2367] = 16'h0000;
initial mem[2368] = 16'h0000;
initial mem[2369] = 16'h0000;
initial mem[2370] = 16'h0000;
initial mem[2371] = 16'h0000;
initial mem[2372] = 16'h0000;
initial mem[2373] = 16'h0000;
initial mem[2374] = 16'h0000;
initial mem[2375] = 16'h0000;
initial mem[2376] = 16'h0000;
initial mem[2377] = 16'h0000;
initial mem[2378] = 16'h0000;
initial mem[2379] = 16'h0000;
initial mem[2380] = 16'h0000;
initial mem[2381] = 16'h0000;
initial mem[2382] = 16'h0000;
initial mem[2383] = 16'h0000;
initial mem[2384] = 16'h0000;
initial mem[2385] = 16'h0000;
initial mem[2386] = 16'h0000;
initial mem[2387] = 16'h0000;
initial mem[2388] = 16'h0000;
initial mem[2389] = 16'h0000;
initial mem[2390] = 16'h0000;
initial mem[2391] = 16'h0000;
initial mem[2392] = 16'h0000;
initial mem[2393] = 16'h0000;
initial mem[2394] = 16'h0000;
initial mem[2395] = 16'h0000;
initial mem[2396] = 16'h0000;
initial mem[2397] = 16'h0000;
initial mem[2398] = 16'h0000;
initial mem[2399] = 16'h0000;
initial mem[2400] = 16'h0000;
initial mem[2401] = 16'h0000;
initial mem[2402] = 16'h0000;
initial mem[2403] = 16'h0000;
initial mem[2404] = 16'h0000;
initial mem[2405] = 16'h0000;
initial mem[2406] = 16'h0000;
initial mem[2407] = 16'h0000;
initial mem[2408] = 16'h0000;
initial mem[2409] = 16'h0000;
initial mem[2410] = 16'h0000;
initial mem[2411] = 16'h0000;
initial mem[2412] = 16'h0000;
initial mem[2413] = 16'h0000;
initial mem[2414] = 16'h0000;
initial mem[2415] = 16'h0000;
initial mem[2416] = 16'h0000;
initial mem[2417] = 16'h0000;
initial mem[2418] = 16'h0000;
initial mem[2419] = 16'h0000;
initial mem[2420] = 16'h0000;
initial mem[2421] = 16'h0000;
initial mem[2422] = 16'h0000;
initial mem[2423] = 16'h0000;
initial mem[2424] = 16'h0000;
initial mem[2425] = 16'h0000;
initial mem[2426] = 16'h0000;
initial mem[2427] = 16'h0000;
initial mem[2428] = 16'h0000;
initial mem[2429] = 16'h0000;
initial mem[2430] = 16'h0000;
initial mem[2431] = 16'h0000;
initial mem[2432] = 16'h0000;
initial mem[2433] = 16'h0000;
initial mem[2434] = 16'h0000;
initial mem[2435] = 16'h0000;
initial mem[2436] = 16'h0000;
initial mem[2437] = 16'h0000;
initial mem[2438] = 16'h0000;
initial mem[2439] = 16'h0000;
initial mem[2440] = 16'h0000;
initial mem[2441] = 16'h0000;
initial mem[2442] = 16'h0000;
initial mem[2443] = 16'h0000;
initial mem[2444] = 16'h0000;
initial mem[2445] = 16'h0000;
initial mem[2446] = 16'h0000;
initial mem[2447] = 16'h0000;
initial mem[2448] = 16'h0000;
initial mem[2449] = 16'h0000;
initial mem[2450] = 16'h0000;
initial mem[2451] = 16'h0000;
initial mem[2452] = 16'h0000;
initial mem[2453] = 16'h0000;
initial mem[2454] = 16'h0000;
initial mem[2455] = 16'h0000;
initial mem[2456] = 16'h0000;
initial mem[2457] = 16'h0000;
initial mem[2458] = 16'h0000;
initial mem[2459] = 16'h0000;
initial mem[2460] = 16'h0000;
initial mem[2461] = 16'h0000;
initial mem[2462] = 16'h0000;
initial mem[2463] = 16'h0000;
initial mem[2464] = 16'h0000;
initial mem[2465] = 16'h0000;
initial mem[2466] = 16'h0000;
initial mem[2467] = 16'h0000;
initial mem[2468] = 16'h0000;
initial mem[2469] = 16'h0000;
initial mem[2470] = 16'h0000;
initial mem[2471] = 16'h0000;
initial mem[2472] = 16'h0000;
initial mem[2473] = 16'h0000;
initial mem[2474] = 16'h0000;
initial mem[2475] = 16'h0000;
initial mem[2476] = 16'h0000;
initial mem[2477] = 16'h0000;
initial mem[2478] = 16'h0000;
initial mem[2479] = 16'h0000;
initial mem[2480] = 16'h0000;
initial mem[2481] = 16'h0000;
initial mem[2482] = 16'h0000;
initial mem[2483] = 16'h0000;
initial mem[2484] = 16'h0000;
initial mem[2485] = 16'h0000;
initial mem[2486] = 16'h0000;
initial mem[2487] = 16'h0000;
initial mem[2488] = 16'h0000;
initial mem[2489] = 16'h0000;
initial mem[2490] = 16'h0000;
initial mem[2491] = 16'h0000;
initial mem[2492] = 16'h0000;
initial mem[2493] = 16'h0000;
initial mem[2494] = 16'h0000;
initial mem[2495] = 16'h0000;
initial mem[2496] = 16'h0000;
initial mem[2497] = 16'h0000;
initial mem[2498] = 16'h0000;
initial mem[2499] = 16'h0000;
initial mem[2500] = 16'h0000;
initial mem[2501] = 16'h0000;
initial mem[2502] = 16'h0000;
initial mem[2503] = 16'h0000;
initial mem[2504] = 16'h0000;
initial mem[2505] = 16'h0000;
initial mem[2506] = 16'h0000;
initial mem[2507] = 16'h0000;
initial mem[2508] = 16'h0000;
initial mem[2509] = 16'h0000;
initial mem[2510] = 16'h0000;
initial mem[2511] = 16'h0000;
initial mem[2512] = 16'h0000;
initial mem[2513] = 16'h0000;
initial mem[2514] = 16'h0000;
initial mem[2515] = 16'h0000;
initial mem[2516] = 16'h0000;
initial mem[2517] = 16'h0000;
initial mem[2518] = 16'h0000;
initial mem[2519] = 16'h0000;
initial mem[2520] = 16'h0000;
initial mem[2521] = 16'h0000;
initial mem[2522] = 16'h0000;
initial mem[2523] = 16'h0000;
initial mem[2524] = 16'h0000;
initial mem[2525] = 16'h0000;
initial mem[2526] = 16'h0000;
initial mem[2527] = 16'h0000;
initial mem[2528] = 16'h0000;
initial mem[2529] = 16'h0000;
initial mem[2530] = 16'h0000;
initial mem[2531] = 16'h0000;
initial mem[2532] = 16'h0000;
initial mem[2533] = 16'h0000;
initial mem[2534] = 16'h0000;
initial mem[2535] = 16'h0000;
initial mem[2536] = 16'h0000;
initial mem[2537] = 16'h0000;
initial mem[2538] = 16'h0000;
initial mem[2539] = 16'h0000;
initial mem[2540] = 16'h0000;
initial mem[2541] = 16'h0000;
initial mem[2542] = 16'h0000;
initial mem[2543] = 16'h0000;
initial mem[2544] = 16'h0000;
initial mem[2545] = 16'h0000;
initial mem[2546] = 16'h0000;
initial mem[2547] = 16'h0000;
initial mem[2548] = 16'h0000;
initial mem[2549] = 16'h0000;
initial mem[2550] = 16'h0000;
initial mem[2551] = 16'h0000;
initial mem[2552] = 16'h0000;
initial mem[2553] = 16'h0000;
initial mem[2554] = 16'h0000;
initial mem[2555] = 16'h0000;
initial mem[2556] = 16'h0000;
initial mem[2557] = 16'h0000;
initial mem[2558] = 16'h0000;
initial mem[2559] = 16'h0000;
initial mem[2560] = 16'h0000;
initial mem[2561] = 16'h0000;
initial mem[2562] = 16'h0000;
initial mem[2563] = 16'h0000;
initial mem[2564] = 16'h0000;
initial mem[2565] = 16'h0000;
initial mem[2566] = 16'h0000;
initial mem[2567] = 16'h0000;
initial mem[2568] = 16'h0000;
initial mem[2569] = 16'h0000;
initial mem[2570] = 16'h0000;
initial mem[2571] = 16'h0000;
initial mem[2572] = 16'h0000;
initial mem[2573] = 16'h0000;
initial mem[2574] = 16'h0000;
initial mem[2575] = 16'h0000;
initial mem[2576] = 16'h0000;
initial mem[2577] = 16'h0000;
initial mem[2578] = 16'h0000;
initial mem[2579] = 16'h0000;
initial mem[2580] = 16'h0000;
initial mem[2581] = 16'h0000;
initial mem[2582] = 16'h0000;
initial mem[2583] = 16'h0000;
initial mem[2584] = 16'h0000;
initial mem[2585] = 16'h0000;
initial mem[2586] = 16'h0000;
initial mem[2587] = 16'h0000;
initial mem[2588] = 16'h0000;
initial mem[2589] = 16'h0000;
initial mem[2590] = 16'h0000;
initial mem[2591] = 16'h0000;
initial mem[2592] = 16'h0000;
initial mem[2593] = 16'h0000;
initial mem[2594] = 16'h0000;
initial mem[2595] = 16'h0000;
initial mem[2596] = 16'h0000;
initial mem[2597] = 16'h0000;
initial mem[2598] = 16'h0000;
initial mem[2599] = 16'h0000;
initial mem[2600] = 16'h0000;
initial mem[2601] = 16'h0000;
initial mem[2602] = 16'h0000;
initial mem[2603] = 16'h0000;
initial mem[2604] = 16'h0000;
initial mem[2605] = 16'h0000;
initial mem[2606] = 16'h0000;
initial mem[2607] = 16'h0000;
initial mem[2608] = 16'h0000;
initial mem[2609] = 16'h0000;
initial mem[2610] = 16'h0000;
initial mem[2611] = 16'h0000;
initial mem[2612] = 16'h0000;
initial mem[2613] = 16'h0000;
initial mem[2614] = 16'h0000;
initial mem[2615] = 16'h0000;
initial mem[2616] = 16'h0000;
initial mem[2617] = 16'h0000;
initial mem[2618] = 16'h0000;
initial mem[2619] = 16'h0000;
initial mem[2620] = 16'h0000;
initial mem[2621] = 16'h0000;
initial mem[2622] = 16'h0000;
initial mem[2623] = 16'h0000;
initial mem[2624] = 16'h0000;
initial mem[2625] = 16'h0000;
initial mem[2626] = 16'h0000;
initial mem[2627] = 16'h0000;
initial mem[2628] = 16'h0000;
initial mem[2629] = 16'h0000;
initial mem[2630] = 16'h0000;
initial mem[2631] = 16'h0000;
initial mem[2632] = 16'h0000;
initial mem[2633] = 16'h0000;
initial mem[2634] = 16'h0000;
initial mem[2635] = 16'h0000;
initial mem[2636] = 16'h0000;
initial mem[2637] = 16'h0000;
initial mem[2638] = 16'h0000;
initial mem[2639] = 16'h0000;
initial mem[2640] = 16'h0000;
initial mem[2641] = 16'h0000;
initial mem[2642] = 16'h0000;
initial mem[2643] = 16'h0000;
initial mem[2644] = 16'h0000;
initial mem[2645] = 16'h0000;
initial mem[2646] = 16'h0000;
initial mem[2647] = 16'h0000;
initial mem[2648] = 16'h0000;
initial mem[2649] = 16'h0000;
initial mem[2650] = 16'h0000;
initial mem[2651] = 16'h0000;
initial mem[2652] = 16'h0000;
initial mem[2653] = 16'h0000;
initial mem[2654] = 16'h0000;
initial mem[2655] = 16'h0000;
initial mem[2656] = 16'h0000;
initial mem[2657] = 16'h0000;
initial mem[2658] = 16'h0000;
initial mem[2659] = 16'h0000;
initial mem[2660] = 16'h0000;
initial mem[2661] = 16'h0000;
initial mem[2662] = 16'h0000;
initial mem[2663] = 16'h0000;
initial mem[2664] = 16'h0000;
initial mem[2665] = 16'h0000;
initial mem[2666] = 16'h0000;
initial mem[2667] = 16'h0000;
initial mem[2668] = 16'h0000;
initial mem[2669] = 16'h0000;
initial mem[2670] = 16'h0000;
initial mem[2671] = 16'h0000;
initial mem[2672] = 16'h0000;
initial mem[2673] = 16'h0000;
initial mem[2674] = 16'h0000;
initial mem[2675] = 16'h0000;
initial mem[2676] = 16'h0000;
initial mem[2677] = 16'h0000;
initial mem[2678] = 16'h0000;
initial mem[2679] = 16'h0000;
initial mem[2680] = 16'h0000;
initial mem[2681] = 16'h0000;
initial mem[2682] = 16'h0000;
initial mem[2683] = 16'h0000;
initial mem[2684] = 16'h0000;
initial mem[2685] = 16'h0000;
initial mem[2686] = 16'h0000;
initial mem[2687] = 16'h0000;
initial mem[2688] = 16'h0000;
initial mem[2689] = 16'h0000;
initial mem[2690] = 16'h0000;
initial mem[2691] = 16'h0000;
initial mem[2692] = 16'h0000;
initial mem[2693] = 16'h0000;
initial mem[2694] = 16'h0000;
initial mem[2695] = 16'h0000;
initial mem[2696] = 16'h0000;
initial mem[2697] = 16'h0000;
initial mem[2698] = 16'h0000;
initial mem[2699] = 16'h0000;
initial mem[2700] = 16'h0000;
initial mem[2701] = 16'h0000;
initial mem[2702] = 16'h0000;
initial mem[2703] = 16'h0000;
initial mem[2704] = 16'h0000;
initial mem[2705] = 16'h0000;
initial mem[2706] = 16'h0000;
initial mem[2707] = 16'h0000;
initial mem[2708] = 16'h0000;
initial mem[2709] = 16'h0000;
initial mem[2710] = 16'h0000;
initial mem[2711] = 16'h0000;
initial mem[2712] = 16'h0000;
initial mem[2713] = 16'h0000;
initial mem[2714] = 16'h0000;
initial mem[2715] = 16'h0000;
initial mem[2716] = 16'h0000;
initial mem[2717] = 16'h0000;
initial mem[2718] = 16'h0000;
initial mem[2719] = 16'h0000;
initial mem[2720] = 16'h0000;
initial mem[2721] = 16'h0000;
initial mem[2722] = 16'h0000;
initial mem[2723] = 16'h0000;
initial mem[2724] = 16'h0000;
initial mem[2725] = 16'h0000;
initial mem[2726] = 16'h0000;
initial mem[2727] = 16'h0000;
initial mem[2728] = 16'h0000;
initial mem[2729] = 16'h0000;
initial mem[2730] = 16'h0000;
initial mem[2731] = 16'h0000;
initial mem[2732] = 16'h0000;
initial mem[2733] = 16'h0000;
initial mem[2734] = 16'h0000;
initial mem[2735] = 16'h0000;
initial mem[2736] = 16'h0000;
initial mem[2737] = 16'h0000;
initial mem[2738] = 16'h0000;
initial mem[2739] = 16'h0000;
initial mem[2740] = 16'h0000;
initial mem[2741] = 16'h0000;
initial mem[2742] = 16'h0000;
initial mem[2743] = 16'h0000;
initial mem[2744] = 16'h0000;
initial mem[2745] = 16'h0000;
initial mem[2746] = 16'h0000;
initial mem[2747] = 16'h0000;
initial mem[2748] = 16'h0000;
initial mem[2749] = 16'h0000;
initial mem[2750] = 16'h0000;
initial mem[2751] = 16'h0000;
initial mem[2752] = 16'h0000;
initial mem[2753] = 16'h0000;
initial mem[2754] = 16'h0000;
initial mem[2755] = 16'h0000;
initial mem[2756] = 16'h0000;
initial mem[2757] = 16'h0000;
initial mem[2758] = 16'h0000;
initial mem[2759] = 16'h0000;
initial mem[2760] = 16'h0000;
initial mem[2761] = 16'h0000;
initial mem[2762] = 16'h0000;
initial mem[2763] = 16'h0000;
initial mem[2764] = 16'h0000;
initial mem[2765] = 16'h0000;
initial mem[2766] = 16'h0000;
initial mem[2767] = 16'h0000;
initial mem[2768] = 16'h0000;
initial mem[2769] = 16'h0000;
initial mem[2770] = 16'h0000;
initial mem[2771] = 16'h0000;
initial mem[2772] = 16'h0000;
initial mem[2773] = 16'h0000;
initial mem[2774] = 16'h0000;
initial mem[2775] = 16'h0000;
initial mem[2776] = 16'h0000;
initial mem[2777] = 16'h0000;
initial mem[2778] = 16'h0000;
initial mem[2779] = 16'h0000;
initial mem[2780] = 16'h0000;
initial mem[2781] = 16'h0000;
initial mem[2782] = 16'h0000;
initial mem[2783] = 16'h0000;
initial mem[2784] = 16'h0000;
initial mem[2785] = 16'h0000;
initial mem[2786] = 16'h0000;
initial mem[2787] = 16'h0000;
initial mem[2788] = 16'h0000;
initial mem[2789] = 16'h0000;
initial mem[2790] = 16'h0000;
initial mem[2791] = 16'h0000;
initial mem[2792] = 16'h0000;
initial mem[2793] = 16'h0000;
initial mem[2794] = 16'h0000;
initial mem[2795] = 16'h0000;
initial mem[2796] = 16'h0000;
initial mem[2797] = 16'h0000;
initial mem[2798] = 16'h0000;
initial mem[2799] = 16'h0000;
initial mem[2800] = 16'h0000;
initial mem[2801] = 16'h0000;
initial mem[2802] = 16'h0000;
initial mem[2803] = 16'h0000;
initial mem[2804] = 16'h0000;
initial mem[2805] = 16'h0000;
initial mem[2806] = 16'h0000;
initial mem[2807] = 16'h0000;
initial mem[2808] = 16'h0000;
initial mem[2809] = 16'h0000;
initial mem[2810] = 16'h0000;
initial mem[2811] = 16'h0000;
initial mem[2812] = 16'h0000;
initial mem[2813] = 16'h0000;
initial mem[2814] = 16'h0000;
initial mem[2815] = 16'h0000;
initial mem[2816] = 16'h0000;
initial mem[2817] = 16'h0000;
initial mem[2818] = 16'h0000;
initial mem[2819] = 16'h0000;
initial mem[2820] = 16'h0000;
initial mem[2821] = 16'h0000;
initial mem[2822] = 16'h0000;
initial mem[2823] = 16'h0000;
initial mem[2824] = 16'h0000;
initial mem[2825] = 16'h0000;
initial mem[2826] = 16'h0000;
initial mem[2827] = 16'h0000;
initial mem[2828] = 16'h0000;
initial mem[2829] = 16'h0000;
initial mem[2830] = 16'h0000;
initial mem[2831] = 16'h0000;
initial mem[2832] = 16'h0000;
initial mem[2833] = 16'h0000;
initial mem[2834] = 16'h0000;
initial mem[2835] = 16'h0000;
initial mem[2836] = 16'h0000;
initial mem[2837] = 16'h0000;
initial mem[2838] = 16'h0000;
initial mem[2839] = 16'h0000;
initial mem[2840] = 16'h0000;
initial mem[2841] = 16'h0000;
initial mem[2842] = 16'h0000;
initial mem[2843] = 16'h0000;
initial mem[2844] = 16'h0000;
initial mem[2845] = 16'h0000;
initial mem[2846] = 16'h0000;
initial mem[2847] = 16'h0000;
initial mem[2848] = 16'h0000;
initial mem[2849] = 16'h0000;
initial mem[2850] = 16'h0000;
initial mem[2851] = 16'h0000;
initial mem[2852] = 16'h0000;
initial mem[2853] = 16'h0000;
initial mem[2854] = 16'h0000;
initial mem[2855] = 16'h0000;
initial mem[2856] = 16'h0000;
initial mem[2857] = 16'h0000;
initial mem[2858] = 16'h0000;
initial mem[2859] = 16'h0000;
initial mem[2860] = 16'h0000;
initial mem[2861] = 16'h0000;
initial mem[2862] = 16'h0000;
initial mem[2863] = 16'h0000;
initial mem[2864] = 16'h0000;
initial mem[2865] = 16'h0000;
initial mem[2866] = 16'h0000;
initial mem[2867] = 16'h0000;
initial mem[2868] = 16'h0000;
initial mem[2869] = 16'h0000;
initial mem[2870] = 16'h0000;
initial mem[2871] = 16'h0000;
initial mem[2872] = 16'h0000;
initial mem[2873] = 16'h0000;
initial mem[2874] = 16'h0000;
initial mem[2875] = 16'h0000;
initial mem[2876] = 16'h0000;
initial mem[2877] = 16'h0000;
initial mem[2878] = 16'h0000;
initial mem[2879] = 16'h0000;
initial mem[2880] = 16'h0000;
initial mem[2881] = 16'h0000;
initial mem[2882] = 16'h0000;
initial mem[2883] = 16'h0000;
initial mem[2884] = 16'h0000;
initial mem[2885] = 16'h0000;
initial mem[2886] = 16'h0000;
initial mem[2887] = 16'h0000;
initial mem[2888] = 16'h0000;
initial mem[2889] = 16'h0000;
initial mem[2890] = 16'h0000;
initial mem[2891] = 16'h0000;
initial mem[2892] = 16'h0000;
initial mem[2893] = 16'h0000;
initial mem[2894] = 16'h0000;
initial mem[2895] = 16'h0000;
initial mem[2896] = 16'h0000;
initial mem[2897] = 16'h0000;
initial mem[2898] = 16'h0000;
initial mem[2899] = 16'h0000;
initial mem[2900] = 16'h0000;
initial mem[2901] = 16'h0000;
initial mem[2902] = 16'h0000;
initial mem[2903] = 16'h0000;
initial mem[2904] = 16'h0000;
initial mem[2905] = 16'h0000;
initial mem[2906] = 16'h0000;
initial mem[2907] = 16'h0000;
initial mem[2908] = 16'h0000;
initial mem[2909] = 16'h0000;
initial mem[2910] = 16'h0000;
initial mem[2911] = 16'h0000;
initial mem[2912] = 16'h0000;
initial mem[2913] = 16'h0000;
initial mem[2914] = 16'h0000;
initial mem[2915] = 16'h0000;
initial mem[2916] = 16'h0000;
initial mem[2917] = 16'h0000;
initial mem[2918] = 16'h0000;
initial mem[2919] = 16'h0000;
initial mem[2920] = 16'h0000;
initial mem[2921] = 16'h0000;
initial mem[2922] = 16'h0000;
initial mem[2923] = 16'h0000;
initial mem[2924] = 16'h0000;
initial mem[2925] = 16'h0000;
initial mem[2926] = 16'h0000;
initial mem[2927] = 16'h0000;
initial mem[2928] = 16'h0000;
initial mem[2929] = 16'h0000;
initial mem[2930] = 16'h0000;
initial mem[2931] = 16'h0000;
initial mem[2932] = 16'h0000;
initial mem[2933] = 16'h0000;
initial mem[2934] = 16'h0000;
initial mem[2935] = 16'h0000;
initial mem[2936] = 16'h0000;
initial mem[2937] = 16'h0000;
initial mem[2938] = 16'h0000;
initial mem[2939] = 16'h0000;
initial mem[2940] = 16'h0000;
initial mem[2941] = 16'h0000;
initial mem[2942] = 16'h0000;
initial mem[2943] = 16'h0000;
initial mem[2944] = 16'h0000;
initial mem[2945] = 16'h0000;
initial mem[2946] = 16'h0000;
initial mem[2947] = 16'h0000;
initial mem[2948] = 16'h0000;
initial mem[2949] = 16'h0000;
initial mem[2950] = 16'h0000;
initial mem[2951] = 16'h0000;
initial mem[2952] = 16'h0000;
initial mem[2953] = 16'h0000;
initial mem[2954] = 16'h0000;
initial mem[2955] = 16'h0000;
initial mem[2956] = 16'h0000;
initial mem[2957] = 16'h0000;
initial mem[2958] = 16'h0000;
initial mem[2959] = 16'h0000;
initial mem[2960] = 16'h0000;
initial mem[2961] = 16'h0000;
initial mem[2962] = 16'h0000;
initial mem[2963] = 16'h0000;
initial mem[2964] = 16'h0000;
initial mem[2965] = 16'h0000;
initial mem[2966] = 16'h0000;
initial mem[2967] = 16'h0000;
initial mem[2968] = 16'h0000;
initial mem[2969] = 16'h0000;
initial mem[2970] = 16'h0000;
initial mem[2971] = 16'h0000;
initial mem[2972] = 16'h0000;
initial mem[2973] = 16'h0000;
initial mem[2974] = 16'h0000;
initial mem[2975] = 16'h0000;
initial mem[2976] = 16'h0000;
initial mem[2977] = 16'h0000;
initial mem[2978] = 16'h0000;
initial mem[2979] = 16'h0000;
initial mem[2980] = 16'h0000;
initial mem[2981] = 16'h0000;
initial mem[2982] = 16'h0000;
initial mem[2983] = 16'h0000;
initial mem[2984] = 16'h0000;
initial mem[2985] = 16'h0000;
initial mem[2986] = 16'h0000;
initial mem[2987] = 16'h0000;
initial mem[2988] = 16'h0000;
initial mem[2989] = 16'h0000;
initial mem[2990] = 16'h0000;
initial mem[2991] = 16'h0000;
initial mem[2992] = 16'h0000;
initial mem[2993] = 16'h0000;
initial mem[2994] = 16'h0000;
initial mem[2995] = 16'h0000;
initial mem[2996] = 16'h0000;
initial mem[2997] = 16'h0000;
initial mem[2998] = 16'h0000;
initial mem[2999] = 16'h0000;
initial mem[3000] = 16'h0000;
initial mem[3001] = 16'h0000;
initial mem[3002] = 16'h0000;
initial mem[3003] = 16'h0000;
initial mem[3004] = 16'h0000;
initial mem[3005] = 16'h0000;
initial mem[3006] = 16'h0000;
initial mem[3007] = 16'h0000;
initial mem[3008] = 16'h0000;
initial mem[3009] = 16'h0000;
initial mem[3010] = 16'h0000;
initial mem[3011] = 16'h0000;
initial mem[3012] = 16'h0000;
initial mem[3013] = 16'h0000;
initial mem[3014] = 16'h0000;
initial mem[3015] = 16'h0000;
initial mem[3016] = 16'h0000;
initial mem[3017] = 16'h0000;
initial mem[3018] = 16'h0000;
initial mem[3019] = 16'h0000;
initial mem[3020] = 16'h0000;
initial mem[3021] = 16'h0000;
initial mem[3022] = 16'h0000;
initial mem[3023] = 16'h0000;
initial mem[3024] = 16'h0000;
initial mem[3025] = 16'h0000;
initial mem[3026] = 16'h0000;
initial mem[3027] = 16'h0000;
initial mem[3028] = 16'h0000;
initial mem[3029] = 16'h0000;
initial mem[3030] = 16'h0000;
initial mem[3031] = 16'h0000;
initial mem[3032] = 16'h0000;
initial mem[3033] = 16'h0000;
initial mem[3034] = 16'h0000;
initial mem[3035] = 16'h0000;
initial mem[3036] = 16'h0000;
initial mem[3037] = 16'h0000;
initial mem[3038] = 16'h0000;
initial mem[3039] = 16'h0000;
initial mem[3040] = 16'h0000;
initial mem[3041] = 16'h0000;
initial mem[3042] = 16'h0000;
initial mem[3043] = 16'h0000;
initial mem[3044] = 16'h0000;
initial mem[3045] = 16'h0000;
initial mem[3046] = 16'h0000;
initial mem[3047] = 16'h0000;
initial mem[3048] = 16'h0000;
initial mem[3049] = 16'h0000;
initial mem[3050] = 16'h0000;
initial mem[3051] = 16'h0000;
initial mem[3052] = 16'h0000;
initial mem[3053] = 16'h0000;
initial mem[3054] = 16'h0000;
initial mem[3055] = 16'h0000;
initial mem[3056] = 16'h0000;
initial mem[3057] = 16'h0000;
initial mem[3058] = 16'h0000;
initial mem[3059] = 16'h0000;
initial mem[3060] = 16'h0000;
initial mem[3061] = 16'h0000;
initial mem[3062] = 16'h0000;
initial mem[3063] = 16'h0000;
initial mem[3064] = 16'h0000;
initial mem[3065] = 16'h0000;
initial mem[3066] = 16'h0000;
initial mem[3067] = 16'h0000;
initial mem[3068] = 16'h0000;
initial mem[3069] = 16'h0000;
initial mem[3070] = 16'h0000;
initial mem[3071] = 16'h0000;
initial mem[3072] = 16'h0000;
initial mem[3073] = 16'h0000;
initial mem[3074] = 16'h0000;
initial mem[3075] = 16'h0000;
initial mem[3076] = 16'h0000;
initial mem[3077] = 16'h0000;
initial mem[3078] = 16'h0000;
initial mem[3079] = 16'h0000;
initial mem[3080] = 16'h0000;
initial mem[3081] = 16'h0000;
initial mem[3082] = 16'h0000;
initial mem[3083] = 16'h0000;
initial mem[3084] = 16'h0000;
initial mem[3085] = 16'h0000;
initial mem[3086] = 16'h0000;
initial mem[3087] = 16'h0000;
initial mem[3088] = 16'h0000;
initial mem[3089] = 16'h0000;
initial mem[3090] = 16'h0000;
initial mem[3091] = 16'h0000;
initial mem[3092] = 16'h0000;
initial mem[3093] = 16'h0000;
initial mem[3094] = 16'h0000;
initial mem[3095] = 16'h0000;
initial mem[3096] = 16'h0000;
initial mem[3097] = 16'h0000;
initial mem[3098] = 16'h0000;
initial mem[3099] = 16'h0000;
initial mem[3100] = 16'h0000;
initial mem[3101] = 16'h0000;
initial mem[3102] = 16'h0000;
initial mem[3103] = 16'h0000;
initial mem[3104] = 16'h0000;
initial mem[3105] = 16'h0000;
initial mem[3106] = 16'h0000;
initial mem[3107] = 16'h0000;
initial mem[3108] = 16'h0000;
initial mem[3109] = 16'h0000;
initial mem[3110] = 16'h0000;
initial mem[3111] = 16'h0000;
initial mem[3112] = 16'h0000;
initial mem[3113] = 16'h0000;
initial mem[3114] = 16'h0000;
initial mem[3115] = 16'h0000;
initial mem[3116] = 16'h0000;
initial mem[3117] = 16'h0000;
initial mem[3118] = 16'h0000;
initial mem[3119] = 16'h0000;
initial mem[3120] = 16'h0000;
initial mem[3121] = 16'h0000;
initial mem[3122] = 16'h0000;
initial mem[3123] = 16'h0000;
initial mem[3124] = 16'h0000;
initial mem[3125] = 16'h0000;
initial mem[3126] = 16'h0000;
initial mem[3127] = 16'h0000;
initial mem[3128] = 16'h0000;
initial mem[3129] = 16'h0000;
initial mem[3130] = 16'h0000;
initial mem[3131] = 16'h0000;
initial mem[3132] = 16'h0000;
initial mem[3133] = 16'h0000;
initial mem[3134] = 16'h0000;
initial mem[3135] = 16'h0000;
initial mem[3136] = 16'h0000;
initial mem[3137] = 16'h0000;
initial mem[3138] = 16'h0000;
initial mem[3139] = 16'h0000;
initial mem[3140] = 16'h0000;
initial mem[3141] = 16'h0000;
initial mem[3142] = 16'h0000;
initial mem[3143] = 16'h0000;
initial mem[3144] = 16'h0000;
initial mem[3145] = 16'h0000;
initial mem[3146] = 16'h0000;
initial mem[3147] = 16'h0000;
initial mem[3148] = 16'h0000;
initial mem[3149] = 16'h0000;
initial mem[3150] = 16'h0000;
initial mem[3151] = 16'h0000;
initial mem[3152] = 16'h0000;
initial mem[3153] = 16'h0000;
initial mem[3154] = 16'h0000;
initial mem[3155] = 16'h0000;
initial mem[3156] = 16'h0000;
initial mem[3157] = 16'h0000;
initial mem[3158] = 16'h0000;
initial mem[3159] = 16'h0000;
initial mem[3160] = 16'h0000;
initial mem[3161] = 16'h0000;
initial mem[3162] = 16'h0000;
initial mem[3163] = 16'h0000;
initial mem[3164] = 16'h0000;
initial mem[3165] = 16'h0000;
initial mem[3166] = 16'h0000;
initial mem[3167] = 16'h0000;
initial mem[3168] = 16'h0000;
initial mem[3169] = 16'h0000;
initial mem[3170] = 16'h0000;
initial mem[3171] = 16'h0000;
initial mem[3172] = 16'h0000;
initial mem[3173] = 16'h0000;
initial mem[3174] = 16'h0000;
initial mem[3175] = 16'h0000;
initial mem[3176] = 16'h0000;
initial mem[3177] = 16'h0000;
initial mem[3178] = 16'h0000;
initial mem[3179] = 16'h0000;
initial mem[3180] = 16'h0000;
initial mem[3181] = 16'h0000;
initial mem[3182] = 16'h0000;
initial mem[3183] = 16'h0000;
initial mem[3184] = 16'h0000;
initial mem[3185] = 16'h0000;
initial mem[3186] = 16'h0000;
initial mem[3187] = 16'h0000;
initial mem[3188] = 16'h0000;
initial mem[3189] = 16'h0000;
initial mem[3190] = 16'h0000;
initial mem[3191] = 16'h0000;
initial mem[3192] = 16'h0000;
initial mem[3193] = 16'h0000;
initial mem[3194] = 16'h0000;
initial mem[3195] = 16'h0000;
initial mem[3196] = 16'h0000;
initial mem[3197] = 16'h0000;
initial mem[3198] = 16'h0000;
initial mem[3199] = 16'h0000;
initial mem[3200] = 16'h0000;
initial mem[3201] = 16'h0000;
initial mem[3202] = 16'h0000;
initial mem[3203] = 16'h0000;
initial mem[3204] = 16'h0000;
initial mem[3205] = 16'h0000;
initial mem[3206] = 16'h0000;
initial mem[3207] = 16'h0000;
initial mem[3208] = 16'h0000;
initial mem[3209] = 16'h0000;
initial mem[3210] = 16'h0000;
initial mem[3211] = 16'h0000;
initial mem[3212] = 16'h0000;
initial mem[3213] = 16'h0000;
initial mem[3214] = 16'h0000;
initial mem[3215] = 16'h0000;
initial mem[3216] = 16'h0000;
initial mem[3217] = 16'h0000;
initial mem[3218] = 16'h0000;
initial mem[3219] = 16'h0000;
initial mem[3220] = 16'h0000;
initial mem[3221] = 16'h0000;
initial mem[3222] = 16'h0000;
initial mem[3223] = 16'h0000;
initial mem[3224] = 16'h0000;
initial mem[3225] = 16'h0000;
initial mem[3226] = 16'h0000;
initial mem[3227] = 16'h0000;
initial mem[3228] = 16'h0000;
initial mem[3229] = 16'h0000;
initial mem[3230] = 16'h0000;
initial mem[3231] = 16'h0000;
initial mem[3232] = 16'h0000;
initial mem[3233] = 16'h0000;
initial mem[3234] = 16'h0000;
initial mem[3235] = 16'h0000;
initial mem[3236] = 16'h0000;
initial mem[3237] = 16'h0000;
initial mem[3238] = 16'h0000;
initial mem[3239] = 16'h0000;
initial mem[3240] = 16'h0000;
initial mem[3241] = 16'h0000;
initial mem[3242] = 16'h0000;
initial mem[3243] = 16'h0000;
initial mem[3244] = 16'h0000;
initial mem[3245] = 16'h0000;
initial mem[3246] = 16'h0000;
initial mem[3247] = 16'h0000;
initial mem[3248] = 16'h0000;
initial mem[3249] = 16'h0000;
initial mem[3250] = 16'h0000;
initial mem[3251] = 16'h0000;
initial mem[3252] = 16'h0000;
initial mem[3253] = 16'h0000;
initial mem[3254] = 16'h0000;
initial mem[3255] = 16'h0000;
initial mem[3256] = 16'h0000;
initial mem[3257] = 16'h0000;
initial mem[3258] = 16'h0000;
initial mem[3259] = 16'h0000;
initial mem[3260] = 16'h0000;
initial mem[3261] = 16'h0000;
initial mem[3262] = 16'h0000;
initial mem[3263] = 16'h0000;
initial mem[3264] = 16'h0000;
initial mem[3265] = 16'h0000;
initial mem[3266] = 16'h0000;
initial mem[3267] = 16'h0000;
initial mem[3268] = 16'h0000;
initial mem[3269] = 16'h0000;
initial mem[3270] = 16'h0000;
initial mem[3271] = 16'h0000;
initial mem[3272] = 16'h0000;
initial mem[3273] = 16'h0000;
initial mem[3274] = 16'h0000;
initial mem[3275] = 16'h0000;
initial mem[3276] = 16'h0000;
initial mem[3277] = 16'h0000;
initial mem[3278] = 16'h0000;
initial mem[3279] = 16'h0000;
initial mem[3280] = 16'h0000;
initial mem[3281] = 16'h0000;
initial mem[3282] = 16'h0000;
initial mem[3283] = 16'h0000;
initial mem[3284] = 16'h0000;
initial mem[3285] = 16'h0000;
initial mem[3286] = 16'h0000;
initial mem[3287] = 16'h0000;
initial mem[3288] = 16'h0000;
initial mem[3289] = 16'h0000;
initial mem[3290] = 16'h0000;
initial mem[3291] = 16'h0000;
initial mem[3292] = 16'h0000;
initial mem[3293] = 16'h0000;
initial mem[3294] = 16'h0000;
initial mem[3295] = 16'h0000;
initial mem[3296] = 16'h0000;
initial mem[3297] = 16'h0000;
initial mem[3298] = 16'h0000;
initial mem[3299] = 16'h0000;
initial mem[3300] = 16'h0000;
initial mem[3301] = 16'h0000;
initial mem[3302] = 16'h0000;
initial mem[3303] = 16'h0000;
initial mem[3304] = 16'h0000;
initial mem[3305] = 16'h0000;
initial mem[3306] = 16'h0000;
initial mem[3307] = 16'h0000;
initial mem[3308] = 16'h0000;
initial mem[3309] = 16'h0000;
initial mem[3310] = 16'h0000;
initial mem[3311] = 16'h0000;
initial mem[3312] = 16'h0000;
initial mem[3313] = 16'h0000;
initial mem[3314] = 16'h0000;
initial mem[3315] = 16'h0000;
initial mem[3316] = 16'h0000;
initial mem[3317] = 16'h0000;
initial mem[3318] = 16'h0000;
initial mem[3319] = 16'h0000;
initial mem[3320] = 16'h0000;
initial mem[3321] = 16'h0000;
initial mem[3322] = 16'h0000;
initial mem[3323] = 16'h0000;
initial mem[3324] = 16'h0000;
initial mem[3325] = 16'h0000;
initial mem[3326] = 16'h0000;
initial mem[3327] = 16'h0000;
initial mem[3328] = 16'h0000;
initial mem[3329] = 16'h0000;
initial mem[3330] = 16'h0000;
initial mem[3331] = 16'h0000;
initial mem[3332] = 16'h0000;
initial mem[3333] = 16'h0000;
initial mem[3334] = 16'h0000;
initial mem[3335] = 16'h0000;
initial mem[3336] = 16'h0000;
initial mem[3337] = 16'h0000;
initial mem[3338] = 16'h0000;
initial mem[3339] = 16'h0000;
initial mem[3340] = 16'h0000;
initial mem[3341] = 16'h0000;
initial mem[3342] = 16'h0000;
initial mem[3343] = 16'h0000;
initial mem[3344] = 16'h0000;
initial mem[3345] = 16'h0000;
initial mem[3346] = 16'h0000;
initial mem[3347] = 16'h0000;
initial mem[3348] = 16'h0000;
initial mem[3349] = 16'h0000;
initial mem[3350] = 16'h0000;
initial mem[3351] = 16'h0000;
initial mem[3352] = 16'h0000;
initial mem[3353] = 16'h0000;
initial mem[3354] = 16'h0000;
initial mem[3355] = 16'h0000;
initial mem[3356] = 16'h0000;
initial mem[3357] = 16'h0000;
initial mem[3358] = 16'h0000;
initial mem[3359] = 16'h0000;
initial mem[3360] = 16'h0000;
initial mem[3361] = 16'h0000;
initial mem[3362] = 16'h0000;
initial mem[3363] = 16'h0000;
initial mem[3364] = 16'h0000;
initial mem[3365] = 16'h0000;
initial mem[3366] = 16'h0000;
initial mem[3367] = 16'h0000;
initial mem[3368] = 16'h0000;
initial mem[3369] = 16'h0000;
initial mem[3370] = 16'h0000;
initial mem[3371] = 16'h0000;
initial mem[3372] = 16'h0000;
initial mem[3373] = 16'h0000;
initial mem[3374] = 16'h0000;
initial mem[3375] = 16'h0000;
initial mem[3376] = 16'h0000;
initial mem[3377] = 16'h0000;
initial mem[3378] = 16'h0000;
initial mem[3379] = 16'h0000;
initial mem[3380] = 16'h0000;
initial mem[3381] = 16'h0000;
initial mem[3382] = 16'h0000;
initial mem[3383] = 16'h0000;
initial mem[3384] = 16'h0000;
initial mem[3385] = 16'h0000;
initial mem[3386] = 16'h0000;
initial mem[3387] = 16'h0000;
initial mem[3388] = 16'h0000;
initial mem[3389] = 16'h0000;
initial mem[3390] = 16'h0000;
initial mem[3391] = 16'h0000;
initial mem[3392] = 16'h0000;
initial mem[3393] = 16'h0000;
initial mem[3394] = 16'h0000;
initial mem[3395] = 16'h0000;
initial mem[3396] = 16'h0000;
initial mem[3397] = 16'h0000;
initial mem[3398] = 16'h0000;
initial mem[3399] = 16'h0000;
initial mem[3400] = 16'h0000;
initial mem[3401] = 16'h0000;
initial mem[3402] = 16'h0000;
initial mem[3403] = 16'h0000;
initial mem[3404] = 16'h0000;
initial mem[3405] = 16'h0000;
initial mem[3406] = 16'h0000;
initial mem[3407] = 16'h0000;
initial mem[3408] = 16'h0000;
initial mem[3409] = 16'h0000;
initial mem[3410] = 16'h0000;
initial mem[3411] = 16'h0000;
initial mem[3412] = 16'h0000;
initial mem[3413] = 16'h0000;
initial mem[3414] = 16'h0000;
initial mem[3415] = 16'h0000;
initial mem[3416] = 16'h0000;
initial mem[3417] = 16'h0000;
initial mem[3418] = 16'h0000;
initial mem[3419] = 16'h0000;
initial mem[3420] = 16'h0000;
initial mem[3421] = 16'h0000;
initial mem[3422] = 16'h0000;
initial mem[3423] = 16'h0000;
initial mem[3424] = 16'h0000;
initial mem[3425] = 16'h0000;
initial mem[3426] = 16'h0000;
initial mem[3427] = 16'h0000;
initial mem[3428] = 16'h0000;
initial mem[3429] = 16'h0000;
initial mem[3430] = 16'h0000;
initial mem[3431] = 16'h0000;
initial mem[3432] = 16'h0000;
initial mem[3433] = 16'h0000;
initial mem[3434] = 16'h0000;
initial mem[3435] = 16'h0000;
initial mem[3436] = 16'h0000;
initial mem[3437] = 16'h0000;
initial mem[3438] = 16'h0000;
initial mem[3439] = 16'h0000;
initial mem[3440] = 16'h0000;
initial mem[3441] = 16'h0000;
initial mem[3442] = 16'h0000;
initial mem[3443] = 16'h0000;
initial mem[3444] = 16'h0000;
initial mem[3445] = 16'h0000;
initial mem[3446] = 16'h0000;
initial mem[3447] = 16'h0000;
initial mem[3448] = 16'h0000;
initial mem[3449] = 16'h0000;
initial mem[3450] = 16'h0000;
initial mem[3451] = 16'h0000;
initial mem[3452] = 16'h0000;
initial mem[3453] = 16'h0000;
initial mem[3454] = 16'h0000;
initial mem[3455] = 16'h0000;
initial mem[3456] = 16'h0000;
initial mem[3457] = 16'h0000;
initial mem[3458] = 16'h0000;
initial mem[3459] = 16'h0000;
initial mem[3460] = 16'h0000;
initial mem[3461] = 16'h0000;
initial mem[3462] = 16'h0000;
initial mem[3463] = 16'h0000;
initial mem[3464] = 16'h0000;
initial mem[3465] = 16'h0000;
initial mem[3466] = 16'h0000;
initial mem[3467] = 16'h0000;
initial mem[3468] = 16'h0000;
initial mem[3469] = 16'h0000;
initial mem[3470] = 16'h0000;
initial mem[3471] = 16'h0000;
initial mem[3472] = 16'h0000;
initial mem[3473] = 16'h0000;
initial mem[3474] = 16'h0000;
initial mem[3475] = 16'h0000;
initial mem[3476] = 16'h0000;
initial mem[3477] = 16'h0000;
initial mem[3478] = 16'h0000;
initial mem[3479] = 16'h0000;
initial mem[3480] = 16'h0000;
initial mem[3481] = 16'h0000;
initial mem[3482] = 16'h0000;
initial mem[3483] = 16'h0000;
initial mem[3484] = 16'h0000;
initial mem[3485] = 16'h0000;
initial mem[3486] = 16'h0000;
initial mem[3487] = 16'h0000;
initial mem[3488] = 16'h0000;
initial mem[3489] = 16'h0000;
initial mem[3490] = 16'h0000;
initial mem[3491] = 16'h0000;
initial mem[3492] = 16'h0000;
initial mem[3493] = 16'h0000;
initial mem[3494] = 16'h0000;
initial mem[3495] = 16'h0000;
initial mem[3496] = 16'h0000;
initial mem[3497] = 16'h0000;
initial mem[3498] = 16'h0000;
initial mem[3499] = 16'h0000;
initial mem[3500] = 16'h0000;
initial mem[3501] = 16'h0000;
initial mem[3502] = 16'h0000;
initial mem[3503] = 16'h0000;
initial mem[3504] = 16'h0000;
initial mem[3505] = 16'h0000;
initial mem[3506] = 16'h0000;
initial mem[3507] = 16'h0000;
initial mem[3508] = 16'h0000;
initial mem[3509] = 16'h0000;
initial mem[3510] = 16'h0000;
initial mem[3511] = 16'h0000;
initial mem[3512] = 16'h0000;
initial mem[3513] = 16'h0000;
initial mem[3514] = 16'h0000;
initial mem[3515] = 16'h0000;
initial mem[3516] = 16'h0000;
initial mem[3517] = 16'h0000;
initial mem[3518] = 16'h0000;
initial mem[3519] = 16'h0000;
initial mem[3520] = 16'h0000;
initial mem[3521] = 16'h0000;
initial mem[3522] = 16'h0000;
initial mem[3523] = 16'h0000;
initial mem[3524] = 16'h0000;
initial mem[3525] = 16'h0000;
initial mem[3526] = 16'h0000;
initial mem[3527] = 16'h0000;
initial mem[3528] = 16'h0000;
initial mem[3529] = 16'h0000;
initial mem[3530] = 16'h0000;
initial mem[3531] = 16'h0000;
initial mem[3532] = 16'h0000;
initial mem[3533] = 16'h0000;
initial mem[3534] = 16'h0000;
initial mem[3535] = 16'h0000;
initial mem[3536] = 16'h0000;
initial mem[3537] = 16'h0000;
initial mem[3538] = 16'h0000;
initial mem[3539] = 16'h0000;
initial mem[3540] = 16'h0000;
initial mem[3541] = 16'h0000;
initial mem[3542] = 16'h0000;
initial mem[3543] = 16'h0000;
initial mem[3544] = 16'h0000;
initial mem[3545] = 16'h0000;
initial mem[3546] = 16'h0000;
initial mem[3547] = 16'h0000;
initial mem[3548] = 16'h0000;
initial mem[3549] = 16'h0000;
initial mem[3550] = 16'h0000;
initial mem[3551] = 16'h0000;
initial mem[3552] = 16'h0000;
initial mem[3553] = 16'h0000;
initial mem[3554] = 16'h0000;
initial mem[3555] = 16'h0000;
initial mem[3556] = 16'h0000;
initial mem[3557] = 16'h0000;
initial mem[3558] = 16'h0000;
initial mem[3559] = 16'h0000;
initial mem[3560] = 16'h0000;
initial mem[3561] = 16'h0000;
initial mem[3562] = 16'h0000;
initial mem[3563] = 16'h0000;
initial mem[3564] = 16'h0000;
initial mem[3565] = 16'h0000;
initial mem[3566] = 16'h0000;
initial mem[3567] = 16'h0000;
initial mem[3568] = 16'h0000;
initial mem[3569] = 16'h0000;
initial mem[3570] = 16'h0000;
initial mem[3571] = 16'h0000;
initial mem[3572] = 16'h0000;
initial mem[3573] = 16'h0000;
initial mem[3574] = 16'h0000;
initial mem[3575] = 16'h0000;
initial mem[3576] = 16'h0000;
initial mem[3577] = 16'h0000;
initial mem[3578] = 16'h0000;
initial mem[3579] = 16'h0000;
initial mem[3580] = 16'h0000;
initial mem[3581] = 16'h0000;
initial mem[3582] = 16'h0000;
initial mem[3583] = 16'h0000;
initial mem[3584] = 16'h0000;
initial mem[3585] = 16'h0000;
initial mem[3586] = 16'h0000;
initial mem[3587] = 16'h0000;
initial mem[3588] = 16'h0000;
initial mem[3589] = 16'h0000;
initial mem[3590] = 16'h0000;
initial mem[3591] = 16'h0000;
initial mem[3592] = 16'h0000;
initial mem[3593] = 16'h0000;
initial mem[3594] = 16'h0000;
initial mem[3595] = 16'h0000;
initial mem[3596] = 16'h0000;
initial mem[3597] = 16'h0000;
initial mem[3598] = 16'h0000;
initial mem[3599] = 16'h0000;
initial mem[3600] = 16'h0000;
initial mem[3601] = 16'h0000;
initial mem[3602] = 16'h0000;
initial mem[3603] = 16'h0000;
initial mem[3604] = 16'h0000;
initial mem[3605] = 16'h0000;
initial mem[3606] = 16'h0000;
initial mem[3607] = 16'h0000;
initial mem[3608] = 16'h0000;
initial mem[3609] = 16'h0000;
initial mem[3610] = 16'h0000;
initial mem[3611] = 16'h0000;
initial mem[3612] = 16'h0000;
initial mem[3613] = 16'h0000;
initial mem[3614] = 16'h0000;
initial mem[3615] = 16'h0000;
initial mem[3616] = 16'h0000;
initial mem[3617] = 16'h0000;
initial mem[3618] = 16'h0000;
initial mem[3619] = 16'h0000;
initial mem[3620] = 16'h0000;
initial mem[3621] = 16'h0000;
initial mem[3622] = 16'h0000;
initial mem[3623] = 16'h0000;
initial mem[3624] = 16'h0000;
initial mem[3625] = 16'h0000;
initial mem[3626] = 16'h0000;
initial mem[3627] = 16'h0000;
initial mem[3628] = 16'h0000;
initial mem[3629] = 16'h0000;
initial mem[3630] = 16'h0000;
initial mem[3631] = 16'h0000;
initial mem[3632] = 16'h0000;
initial mem[3633] = 16'h0000;
initial mem[3634] = 16'h0000;
initial mem[3635] = 16'h0000;
initial mem[3636] = 16'h0000;
initial mem[3637] = 16'h0000;
initial mem[3638] = 16'h0000;
initial mem[3639] = 16'h0000;
initial mem[3640] = 16'h0000;
initial mem[3641] = 16'h0000;
initial mem[3642] = 16'h0000;
initial mem[3643] = 16'h0000;
initial mem[3644] = 16'h0000;
initial mem[3645] = 16'h0000;
initial mem[3646] = 16'h0000;
initial mem[3647] = 16'h0000;
initial mem[3648] = 16'h0000;
initial mem[3649] = 16'h0000;
initial mem[3650] = 16'h0000;
initial mem[3651] = 16'h0000;
initial mem[3652] = 16'h0000;
initial mem[3653] = 16'h0000;
initial mem[3654] = 16'h0000;
initial mem[3655] = 16'h0000;
initial mem[3656] = 16'h0000;
initial mem[3657] = 16'h0000;
initial mem[3658] = 16'h0000;
initial mem[3659] = 16'h0000;
initial mem[3660] = 16'h0000;
initial mem[3661] = 16'h0000;
initial mem[3662] = 16'h0000;
initial mem[3663] = 16'h0000;
initial mem[3664] = 16'h0000;
initial mem[3665] = 16'h0000;
initial mem[3666] = 16'h0000;
initial mem[3667] = 16'h0000;
initial mem[3668] = 16'h0000;
initial mem[3669] = 16'h0000;
initial mem[3670] = 16'h0000;
initial mem[3671] = 16'h0000;
initial mem[3672] = 16'h0000;
initial mem[3673] = 16'h0000;
initial mem[3674] = 16'h0000;
initial mem[3675] = 16'h0000;
initial mem[3676] = 16'h0000;
initial mem[3677] = 16'h0000;
initial mem[3678] = 16'h0000;
initial mem[3679] = 16'h0000;
initial mem[3680] = 16'h0000;
initial mem[3681] = 16'h0000;
initial mem[3682] = 16'h0000;
initial mem[3683] = 16'h0000;
initial mem[3684] = 16'h0000;
initial mem[3685] = 16'h0000;
initial mem[3686] = 16'h0000;
initial mem[3687] = 16'h0000;
initial mem[3688] = 16'h0000;
initial mem[3689] = 16'h0000;
initial mem[3690] = 16'h0000;
initial mem[3691] = 16'h0000;
initial mem[3692] = 16'h0000;
initial mem[3693] = 16'h0000;
initial mem[3694] = 16'h0000;
initial mem[3695] = 16'h0000;
initial mem[3696] = 16'h0000;
initial mem[3697] = 16'h0000;
initial mem[3698] = 16'h0000;
initial mem[3699] = 16'h0000;
initial mem[3700] = 16'h0000;
initial mem[3701] = 16'h0000;
initial mem[3702] = 16'h0000;
initial mem[3703] = 16'h0000;
initial mem[3704] = 16'h0000;
initial mem[3705] = 16'h0000;
initial mem[3706] = 16'h0000;
initial mem[3707] = 16'h0000;
initial mem[3708] = 16'h0000;
initial mem[3709] = 16'h0000;
initial mem[3710] = 16'h0000;
initial mem[3711] = 16'h0000;
initial mem[3712] = 16'h0000;
initial mem[3713] = 16'h0000;
initial mem[3714] = 16'h0000;
initial mem[3715] = 16'h0000;
initial mem[3716] = 16'h0000;
initial mem[3717] = 16'h0000;
initial mem[3718] = 16'h0000;
initial mem[3719] = 16'h0000;
initial mem[3720] = 16'h0000;
initial mem[3721] = 16'h0000;
initial mem[3722] = 16'h0000;
initial mem[3723] = 16'h0000;
initial mem[3724] = 16'h0000;
initial mem[3725] = 16'h0000;
initial mem[3726] = 16'h0000;
initial mem[3727] = 16'h0000;
initial mem[3728] = 16'h0000;
initial mem[3729] = 16'h0000;
initial mem[3730] = 16'h0000;
initial mem[3731] = 16'h0000;
initial mem[3732] = 16'h0000;
initial mem[3733] = 16'h0000;
initial mem[3734] = 16'h0000;
initial mem[3735] = 16'h0000;
initial mem[3736] = 16'h0000;
initial mem[3737] = 16'h0000;
initial mem[3738] = 16'h0000;
initial mem[3739] = 16'h0000;
initial mem[3740] = 16'h0000;
initial mem[3741] = 16'h0000;
initial mem[3742] = 16'h0000;
initial mem[3743] = 16'h0000;
initial mem[3744] = 16'h0000;
initial mem[3745] = 16'h0000;
initial mem[3746] = 16'h0000;
initial mem[3747] = 16'h0000;
initial mem[3748] = 16'h0000;
initial mem[3749] = 16'h0000;
initial mem[3750] = 16'h0000;
initial mem[3751] = 16'h0000;
initial mem[3752] = 16'h0000;
initial mem[3753] = 16'h0000;
initial mem[3754] = 16'h0000;
initial mem[3755] = 16'h0000;
initial mem[3756] = 16'h0000;
initial mem[3757] = 16'h0000;
initial mem[3758] = 16'h0000;
initial mem[3759] = 16'h0000;
initial mem[3760] = 16'h0000;
initial mem[3761] = 16'h0000;
initial mem[3762] = 16'h0000;
initial mem[3763] = 16'h0000;
initial mem[3764] = 16'h0000;
initial mem[3765] = 16'h0000;
initial mem[3766] = 16'h0000;
initial mem[3767] = 16'h0000;
initial mem[3768] = 16'h0000;
initial mem[3769] = 16'h0000;
initial mem[3770] = 16'h0000;
initial mem[3771] = 16'h0000;
initial mem[3772] = 16'h0000;
initial mem[3773] = 16'h0000;
initial mem[3774] = 16'h0000;
initial mem[3775] = 16'h0000;
initial mem[3776] = 16'h0000;
initial mem[3777] = 16'h0000;
initial mem[3778] = 16'h0000;
initial mem[3779] = 16'h0000;
initial mem[3780] = 16'h0000;
initial mem[3781] = 16'h0000;
initial mem[3782] = 16'h0000;
initial mem[3783] = 16'h0000;
initial mem[3784] = 16'h0000;
initial mem[3785] = 16'h0000;
initial mem[3786] = 16'h0000;
initial mem[3787] = 16'h0000;
initial mem[3788] = 16'h0000;
initial mem[3789] = 16'h0000;
initial mem[3790] = 16'h0000;
initial mem[3791] = 16'h0000;
initial mem[3792] = 16'h0000;
initial mem[3793] = 16'h0000;
initial mem[3794] = 16'h0000;
initial mem[3795] = 16'h0000;
initial mem[3796] = 16'h0000;
initial mem[3797] = 16'h0000;
initial mem[3798] = 16'h0000;
initial mem[3799] = 16'h0000;
initial mem[3800] = 16'h0000;
initial mem[3801] = 16'h0000;
initial mem[3802] = 16'h0000;
initial mem[3803] = 16'h0000;
initial mem[3804] = 16'h0000;
initial mem[3805] = 16'h0000;
initial mem[3806] = 16'h0000;
initial mem[3807] = 16'h0000;
initial mem[3808] = 16'h0000;
initial mem[3809] = 16'h0000;
initial mem[3810] = 16'h0000;
initial mem[3811] = 16'h0000;
initial mem[3812] = 16'h0000;
initial mem[3813] = 16'h0000;
initial mem[3814] = 16'h0000;
initial mem[3815] = 16'h0000;
initial mem[3816] = 16'h0000;
initial mem[3817] = 16'h0000;
initial mem[3818] = 16'h0000;
initial mem[3819] = 16'h0000;
initial mem[3820] = 16'h0000;
initial mem[3821] = 16'h0000;
initial mem[3822] = 16'h0000;
initial mem[3823] = 16'h0000;
initial mem[3824] = 16'h0000;
initial mem[3825] = 16'h0000;
initial mem[3826] = 16'h0000;
initial mem[3827] = 16'h0000;
initial mem[3828] = 16'h0000;
initial mem[3829] = 16'h0000;
initial mem[3830] = 16'h0000;
initial mem[3831] = 16'h0000;
initial mem[3832] = 16'h0000;
initial mem[3833] = 16'h0000;
initial mem[3834] = 16'h0000;
initial mem[3835] = 16'h0000;
initial mem[3836] = 16'h0000;
initial mem[3837] = 16'h0000;
initial mem[3838] = 16'h0000;
initial mem[3839] = 16'h0000;
initial mem[3840] = 16'h0000;
initial mem[3841] = 16'h0000;
initial mem[3842] = 16'h0000;
initial mem[3843] = 16'h0000;
initial mem[3844] = 16'h0000;
initial mem[3845] = 16'h0000;
initial mem[3846] = 16'h0000;
initial mem[3847] = 16'h0000;
initial mem[3848] = 16'h0000;
initial mem[3849] = 16'h0000;
initial mem[3850] = 16'h0000;
initial mem[3851] = 16'h0000;
initial mem[3852] = 16'h0000;
initial mem[3853] = 16'h0000;
initial mem[3854] = 16'h0000;
initial mem[3855] = 16'h0000;
initial mem[3856] = 16'h0000;
initial mem[3857] = 16'h0000;
initial mem[3858] = 16'h0000;
initial mem[3859] = 16'h0000;
initial mem[3860] = 16'h0000;
initial mem[3861] = 16'h0000;
initial mem[3862] = 16'h0000;
initial mem[3863] = 16'h0000;
initial mem[3864] = 16'h0000;
initial mem[3865] = 16'h0000;
initial mem[3866] = 16'h0000;
initial mem[3867] = 16'h0000;
initial mem[3868] = 16'h0000;
initial mem[3869] = 16'h0000;
initial mem[3870] = 16'h0000;
initial mem[3871] = 16'h0000;
initial mem[3872] = 16'h0000;
initial mem[3873] = 16'h0000;
initial mem[3874] = 16'h0000;
initial mem[3875] = 16'h0000;
initial mem[3876] = 16'h0000;
initial mem[3877] = 16'h0000;
initial mem[3878] = 16'h0000;
initial mem[3879] = 16'h0000;
initial mem[3880] = 16'h0000;
initial mem[3881] = 16'h0000;
initial mem[3882] = 16'h0000;
initial mem[3883] = 16'h0000;
initial mem[3884] = 16'h0000;
initial mem[3885] = 16'h0000;
initial mem[3886] = 16'h0000;
initial mem[3887] = 16'h0000;
initial mem[3888] = 16'h0000;
initial mem[3889] = 16'h0000;
initial mem[3890] = 16'h0000;
initial mem[3891] = 16'h0000;
initial mem[3892] = 16'h0000;
initial mem[3893] = 16'h0000;
initial mem[3894] = 16'h0000;
initial mem[3895] = 16'h0000;
initial mem[3896] = 16'h0000;
initial mem[3897] = 16'h0000;
initial mem[3898] = 16'h0000;
initial mem[3899] = 16'h0000;
initial mem[3900] = 16'h0000;
initial mem[3901] = 16'h0000;
initial mem[3902] = 16'h0000;
initial mem[3903] = 16'h0000;
initial mem[3904] = 16'h0000;
initial mem[3905] = 16'h0000;
initial mem[3906] = 16'h0000;
initial mem[3907] = 16'h0000;
initial mem[3908] = 16'h0000;
initial mem[3909] = 16'h0000;
initial mem[3910] = 16'h0000;
initial mem[3911] = 16'h0000;
initial mem[3912] = 16'h0000;
initial mem[3913] = 16'h0000;
initial mem[3914] = 16'h0000;
initial mem[3915] = 16'h0000;
initial mem[3916] = 16'h0000;
initial mem[3917] = 16'h0000;
initial mem[3918] = 16'h0000;
initial mem[3919] = 16'h0000;
initial mem[3920] = 16'h0000;
initial mem[3921] = 16'h0000;
initial mem[3922] = 16'h0000;
initial mem[3923] = 16'h0000;
initial mem[3924] = 16'h0000;
initial mem[3925] = 16'h0000;
initial mem[3926] = 16'h0000;
initial mem[3927] = 16'h0000;
initial mem[3928] = 16'h0000;
initial mem[3929] = 16'h0000;
initial mem[3930] = 16'h0000;
initial mem[3931] = 16'h0000;
initial mem[3932] = 16'h0000;
initial mem[3933] = 16'h0000;
initial mem[3934] = 16'h0000;
initial mem[3935] = 16'h0000;
initial mem[3936] = 16'h0000;
initial mem[3937] = 16'h0000;
initial mem[3938] = 16'h0000;
initial mem[3939] = 16'h0000;
initial mem[3940] = 16'h0000;
initial mem[3941] = 16'h0000;
initial mem[3942] = 16'h0000;
initial mem[3943] = 16'h0000;
initial mem[3944] = 16'h0000;
initial mem[3945] = 16'h0000;
initial mem[3946] = 16'h0000;
initial mem[3947] = 16'h0000;
initial mem[3948] = 16'h0000;
initial mem[3949] = 16'h0000;
initial mem[3950] = 16'h0000;
initial mem[3951] = 16'h0000;
initial mem[3952] = 16'h0000;
initial mem[3953] = 16'h0000;
initial mem[3954] = 16'h0000;
initial mem[3955] = 16'h0000;
initial mem[3956] = 16'h0000;
initial mem[3957] = 16'h0000;
initial mem[3958] = 16'h0000;
initial mem[3959] = 16'h0000;
initial mem[3960] = 16'h0000;
initial mem[3961] = 16'h0000;
initial mem[3962] = 16'h0000;
initial mem[3963] = 16'h0000;
initial mem[3964] = 16'h0000;
initial mem[3965] = 16'h0000;
initial mem[3966] = 16'h0000;
initial mem[3967] = 16'h0000;
initial mem[3968] = 16'h0000;
initial mem[3969] = 16'h0000;
initial mem[3970] = 16'h0000;
initial mem[3971] = 16'h0000;
initial mem[3972] = 16'h0000;
initial mem[3973] = 16'h0000;
initial mem[3974] = 16'h0000;
initial mem[3975] = 16'h0000;
initial mem[3976] = 16'h0000;
initial mem[3977] = 16'h0000;
initial mem[3978] = 16'h0000;
initial mem[3979] = 16'h0000;
initial mem[3980] = 16'h0000;
initial mem[3981] = 16'h0000;
initial mem[3982] = 16'h0000;
initial mem[3983] = 16'h0000;
initial mem[3984] = 16'h0000;
initial mem[3985] = 16'h0000;
initial mem[3986] = 16'h0000;
initial mem[3987] = 16'h0000;
initial mem[3988] = 16'h0000;
initial mem[3989] = 16'h0000;
initial mem[3990] = 16'h0000;
initial mem[3991] = 16'h0000;
initial mem[3992] = 16'h0000;
initial mem[3993] = 16'h0000;
initial mem[3994] = 16'h0000;
initial mem[3995] = 16'h0000;
initial mem[3996] = 16'h0000;
initial mem[3997] = 16'h0000;
initial mem[3998] = 16'h0000;
initial mem[3999] = 16'h0000;
initial mem[4000] = 16'h0000;
initial mem[4001] = 16'h0000;
initial mem[4002] = 16'h0000;
initial mem[4003] = 16'h0000;
initial mem[4004] = 16'h0000;
initial mem[4005] = 16'h0000;
initial mem[4006] = 16'h0000;
initial mem[4007] = 16'h0000;
initial mem[4008] = 16'h0000;
initial mem[4009] = 16'h0000;
initial mem[4010] = 16'h0000;
initial mem[4011] = 16'h0000;
initial mem[4012] = 16'h0000;
initial mem[4013] = 16'h0000;
initial mem[4014] = 16'h0000;
initial mem[4015] = 16'h0000;
initial mem[4016] = 16'h0000;
initial mem[4017] = 16'h0000;
initial mem[4018] = 16'h0000;
initial mem[4019] = 16'h0000;
initial mem[4020] = 16'h0000;
initial mem[4021] = 16'h0000;
initial mem[4022] = 16'h0000;
initial mem[4023] = 16'h0000;
initial mem[4024] = 16'h0000;
initial mem[4025] = 16'h0000;
initial mem[4026] = 16'h0000;
initial mem[4027] = 16'h0000;
initial mem[4028] = 16'h0000;
initial mem[4029] = 16'h0000;
initial mem[4030] = 16'h0000;
initial mem[4031] = 16'h0000;
initial mem[4032] = 16'h0000;
initial mem[4033] = 16'h0000;
initial mem[4034] = 16'h0000;
initial mem[4035] = 16'h0000;
initial mem[4036] = 16'h0000;
initial mem[4037] = 16'h0000;
initial mem[4038] = 16'h0000;
initial mem[4039] = 16'h0000;
initial mem[4040] = 16'h0000;
initial mem[4041] = 16'h0000;
initial mem[4042] = 16'h0000;
initial mem[4043] = 16'h0000;
initial mem[4044] = 16'h0000;
initial mem[4045] = 16'h0000;
initial mem[4046] = 16'h0000;
initial mem[4047] = 16'h0000;
initial mem[4048] = 16'h0000;
initial mem[4049] = 16'h0000;
initial mem[4050] = 16'h0000;
initial mem[4051] = 16'h0000;
initial mem[4052] = 16'h0000;
initial mem[4053] = 16'h0000;
initial mem[4054] = 16'h0000;
initial mem[4055] = 16'h0000;
initial mem[4056] = 16'h0000;
initial mem[4057] = 16'h0000;
initial mem[4058] = 16'h0000;
initial mem[4059] = 16'h0000;
initial mem[4060] = 16'h0000;
initial mem[4061] = 16'h0000;
initial mem[4062] = 16'h0000;
initial mem[4063] = 16'h0000;
initial mem[4064] = 16'h0000;
initial mem[4065] = 16'h0000;
initial mem[4066] = 16'h0000;
initial mem[4067] = 16'h0000;
initial mem[4068] = 16'h0000;
initial mem[4069] = 16'h0000;
initial mem[4070] = 16'h0000;
initial mem[4071] = 16'h0000;
initial mem[4072] = 16'h0000;
initial mem[4073] = 16'h0000;
initial mem[4074] = 16'h0000;
initial mem[4075] = 16'h0000;
initial mem[4076] = 16'h0000;
initial mem[4077] = 16'h0000;
initial mem[4078] = 16'h0000;
initial mem[4079] = 16'h0000;
initial mem[4080] = 16'h0000;
initial mem[4081] = 16'h0000;
initial mem[4082] = 16'h0000;
initial mem[4083] = 16'h0000;
initial mem[4084] = 16'h0000;
initial mem[4085] = 16'h0000;
initial mem[4086] = 16'h0000;
initial mem[4087] = 16'h0000;
initial mem[4088] = 16'h0000;
initial mem[4089] = 16'h0000;
initial mem[4090] = 16'h0000;
initial mem[4091] = 16'h0000;
initial mem[4092] = 16'h0000;
initial mem[4093] = 16'h0000;
initial mem[4094] = 16'h0000;
initial mem[4095] = 16'h0000;
always @(posedge CLK)
begin
       dout <= mem[ADDRESS];
end
endmodule
