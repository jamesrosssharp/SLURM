/*
 *	multiplier placeholder
 *
 *
 */

module mult (
	input [15:0] A,
	input [15:0] B,
	output [31:0] out
);

assign out = A*B;

endmodule
