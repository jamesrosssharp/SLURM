/* boot_memory.v : boot memory */

module boot_memory
#(parameter BITS = 16, ADDRESS_BITS = 8)
(
  input CLK,
  input [ADDRESS_BITS - 1 : 0]  ADDRESS,
  input [BITS - 1 : 0] DATA_IN,
  output [BITS - 1 : 0] DATA_OUT,
  input WR
);

localparam ROM_ADDRESS_BITS = 8;

reg [BITS - 1:0] mem [(1 << ROM_ADDRESS_BITS) - 1:0];
reg [BITS - 1:0] dout;
assign DATA_OUT = dout;
initial mem[0] = 16'h1004;
initial mem[1] = 16'h4e00;
initial mem[2] = 16'h100e;
initial mem[3] = 16'h4e0a;
initial mem[4] = 16'h100e;
initial mem[5] = 16'h4e0a;
initial mem[6] = 16'h100e;
initial mem[7] = 16'h4e0a;
initial mem[8] = 16'h100e;
initial mem[9] = 16'h4e0a;
initial mem[10] = 16'h100e;
initial mem[11] = 16'h4e0a;
initial mem[12] = 16'h0000;
initial mem[13] = 16'h0000;
initial mem[14] = 16'h0000;
initial mem[15] = 16'h0000;
initial mem[16] = 16'h0000;
initial mem[17] = 16'h0000;
initial mem[18] = 16'h0000;
initial mem[19] = 16'h0000;
initial mem[20] = 16'h0000;
initial mem[21] = 16'h0000;
initial mem[22] = 16'h0000;
initial mem[23] = 16'h0000;
initial mem[24] = 16'h0000;
initial mem[25] = 16'h0000;
initial mem[26] = 16'h0000;
initial mem[27] = 16'h0000;
initial mem[28] = 16'h0000;
initial mem[29] = 16'h0000;
initial mem[30] = 16'h0000;
initial mem[31] = 16'h0000;
initial mem[32] = 16'h1002;
initial mem[33] = 16'h3011;
initial mem[34] = 16'hf010;
initial mem[35] = 16'h3012;
initial mem[36] = 16'h1400;
initial mem[37] = 16'hf012;
initial mem[38] = 16'h1002;
initial mem[39] = 16'h3048;
initial mem[40] = 16'h1fff;
initial mem[41] = 16'h303f;
initial mem[42] = 16'h3331;
initial mem[43] = 16'h1005;
initial mem[44] = 16'h4104;
initial mem[45] = 16'h3341;
initial mem[46] = 16'h1005;
initial mem[47] = 16'h4100;
initial mem[48] = 16'h3018;
initial mem[49] = 16'h1400;
initial mem[50] = 16'hf000;
initial mem[51] = 16'h1400;
initial mem[52] = 16'hf011;
initial mem[53] = 16'h1010;
initial mem[54] = 16'h3030;
initial mem[55] = 16'h1400;
initial mem[56] = 16'hf035;
initial mem[57] = 16'h1ff0;
initial mem[58] = 16'h3030;
initial mem[59] = 16'h1400;
initial mem[60] = 16'hf036;
initial mem[61] = 16'h3018;
initial mem[62] = 16'h1700;
initial mem[63] = 16'hf010;
initial mem[64] = 16'h1fff;
initial mem[65] = 16'h309f;
initial mem[66] = 16'h1700;
initial mem[67] = 16'hf091;
initial mem[68] = 16'h0000;
initial mem[69] = 16'h0000;
initial mem[70] = 16'h0000;
initial mem[71] = 16'h0601;
initial mem[72] = 16'h3031;
initial mem[73] = 16'h1400;
initial mem[74] = 16'hf032;
initial mem[75] = 16'h0700;
initial mem[76] = 16'h0000;
initial mem[77] = 16'h0000;
initial mem[78] = 16'h0000;
initial mem[79] = 16'h0000;
initial mem[80] = 16'h0600;
initial mem[81] = 16'h1003;
initial mem[82] = 16'h301f;
initial mem[83] = 16'hf010;
initial mem[84] = 16'h1002;
initial mem[85] = 16'h3048;
initial mem[86] = 16'h1004;
initial mem[87] = 16'h3030;
initial mem[88] = 16'h3331;
initial mem[89] = 16'h100b;
initial mem[90] = 16'h4100;
initial mem[91] = 16'h3341;
initial mem[92] = 16'h100a;
initial mem[93] = 16'h410c;
initial mem[94] = 16'h1400;
initial mem[95] = 16'he014;
initial mem[96] = 16'h2611;
initial mem[97] = 16'h100a;
initial mem[98] = 16'h4002;
initial mem[99] = 16'h1002;
initial mem[100] = 16'h3013;
initial mem[101] = 16'hf010;
initial mem[102] = 16'h1020;
initial mem[103] = 16'h3030;
initial mem[104] = 16'h1020;
initial mem[105] = 16'h3040;
initial mem[106] = 16'ha310;
initial mem[107] = 16'h1010;
initial mem[108] = 16'h4f00;
initial mem[109] = 16'h3131;
initial mem[110] = 16'h3341;
initial mem[111] = 16'h100d;
initial mem[112] = 16'h4104;
initial mem[113] = 16'h1700;
initial mem[114] = 16'hf000;
initial mem[115] = 16'h1020;
initial mem[116] = 16'h4e00;
initial mem[117] = 16'h1400;
initial mem[118] = 16'he084;
initial mem[119] = 16'h1004;
initial mem[120] = 16'h3181;
initial mem[121] = 16'h1000;
initial mem[122] = 16'hf080;
initial mem[123] = 16'h1fff;
initial mem[124] = 16'h309f;
initial mem[125] = 16'h1700;
initial mem[126] = 16'hf091;
initial mem[127] = 16'h0101;
initial mem[128] = 16'h207f;
initial mem[129] = 16'h2041;
initial mem[130] = 16'h0411;
initial mem[131] = 16'h0411;
initial mem[132] = 16'h0411;
initial mem[133] = 16'h0411;
initial mem[134] = 16'h351f;
initial mem[135] = 16'h1012;
initial mem[136] = 16'h4f00;
initial mem[137] = 16'h0000;
initial mem[138] = 16'h2014;
initial mem[139] = 16'h351f;
initial mem[140] = 16'h1012;
initial mem[141] = 16'h4f00;
initial mem[142] = 16'h20f7;
initial mem[143] = 16'h0100;
initial mem[144] = 16'h3c1a;
initial mem[145] = 16'h1012;
initial mem[146] = 16'h420e;
initial mem[147] = 16'h1005;
initial mem[148] = 16'h3117;
initial mem[149] = 16'h1013;
initial mem[150] = 16'h4e02;
initial mem[151] = 16'h1003;
initial mem[152] = 16'h3110;
initial mem[153] = 16'h1000;
initial mem[154] = 16'hf010;
initial mem[155] = 16'h1000;
initial mem[156] = 16'he021;
initial mem[157] = 16'h3d21;
initial mem[158] = 16'h1013;
initial mem[159] = 16'h4006;
initial mem[160] = 16'h0100;
initial mem[161] = 16'h0000;
always @(posedge CLK)
begin
  if (WR == 1'b1) mem[ADDRESS] <= DATA_IN; 
       dout <= mem[ADDRESS];
end
endmodule
